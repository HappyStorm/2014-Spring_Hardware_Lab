`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:13:49 06/22/2014 
// Design Name: 
// Module Name:    LCD_DISPLAY 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module LCD_DISPLAY(LEFT_GRAPH, RIGHT_GRAPH, LCD_CLK, RESETN, LCD_DATA, LCD_ENABLE, LCD_RW, LCD_RSTN, LCD_CS1, LCD_CS2, LCD_DI);
/******************************
 * I/O Port Declare   		   *
 ******************************/
	input [0:4095] LEFT_GRAPH;
	input [0:4095] RIGHT_GRAPH;
	input LCD_CLK;
	input RESETN;
	output reg [7:0]  LCD_DATA;
	output LCD_ENABLE; 
	output reg LCD_RW;
	output LCD_RSTN;
	output reg LCD_CS1 = 1;
	output reg LCD_CS2 = 1;
	output reg LCD_DI;
/******************************
 * Net Declare       		   *
 ******************************/
	reg [7:0]  LCD_DATA_NEXT;
	reg LCD_RW_NEXT;
	reg LCD_DI_NEXT;
	
	reg [2:0] STATE, STATE_NEXT;
	reg [2:0] X_PAGE, X_PAGE_NEXT;
	reg [5:0] Y, Y_NEXT;
	reg [1:0] IMAGE;
	reg [1:0] IMAGE_NEXT;
	reg [7:0] PATTERN;
	reg [8:0]  INDEX, INDEX_NEXT;
	reg [15:0] PAUSE_TIME, PAUSE_TIME_NEXT;
	
	reg START, START_NEXT;	
	reg NEW_PAGE, NEW_PAGE_NEXT;
	reg NEW_COL, NEW_COL_NEXT;
	reg [2:0] PAGE_COUNTER, PAGE_COUNTER_NEXT;
	reg [6:0] COL_COUNTER, COL_COUNTER_NEXT;
	reg ENABLE, ENABLE_NEXT;
	
	//added
	reg LCD_CS1_NEXT, LCD_CS2_NEXT, LCD_SELECT, LCD_SELECT_NEXT, LCD_SIDE, LCD_SIDE_NEXT;
	
	parameter Init = 3'd0, Set_StartLine = 3'd1, Clear_Screen = 3'd2, Copy_Image = 3'd3, Pause = 3'd4;
	parameter Delay = 16'b1000_0000_0000_0000;
	
/******************************
 * Declare   	         	   *
 ******************************/
	assign LCD_ENABLE = LCD_CLK & ENABLE; // when ENABLE=1, LCD write can occur at falling edge of clock
	assign LCD_RSTN = RESETN;
	assign PAUSED_TO_THE_END = (PAUSE_TIME == 0) ? 1 : 0;	
	
	always@(posedge LCD_CLK or negedge RESETN) begin
		if (!RESETN) begin
			STATE    <= Init;
			PAUSE_TIME    <= Delay;
			X_PAGE   <= 0;
			Y  <= 0;
			INDEX 	<=  0;
			LCD_DI   <= 0;
			LCD_RW   <= 0;
			IMAGE    <= 0;
			START <= 0;
			NEW_PAGE <= 1'b0;
			NEW_COL <= 1'b0;
			COL_COUNTER <= 0;
			PAGE_COUNTER <= 0;
			ENABLE <= 1'b0;
			//added
			LCD_CS1 <= 1;
			LCD_CS2 <= 1;
			LCD_SELECT <= 0;
			LCD_SIDE <= 0;
			//added
		end else begin
			STATE    <= STATE_NEXT;
			PAUSE_TIME    <= PAUSE_TIME_NEXT;
			X_PAGE   <= X_PAGE_NEXT;
			Y  <= Y_NEXT;
			INDEX<= INDEX_NEXT;
			LCD_DI   <= LCD_DI_NEXT;
			LCD_RW   <= LCD_RW_NEXT;
			LCD_DATA <= LCD_DATA_NEXT;
			IMAGE <= IMAGE_NEXT;	
			START <= START_NEXT;	
			NEW_PAGE <= NEW_PAGE_NEXT;
			NEW_COL <= NEW_COL_NEXT;
			COL_COUNTER <= COL_COUNTER_NEXT;
			PAGE_COUNTER <= PAGE_COUNTER_NEXT;
			ENABLE <= ENABLE_NEXT;
			//added
			LCD_CS1 <= LCD_CS1_NEXT;
			LCD_CS2 <= LCD_CS2_NEXT;
			LCD_SELECT <= LCD_SELECT_NEXT;
			LCD_SIDE <= LCD_SIDE_NEXT;
			//added
		end
	end

	always @(*) begin
		// default assignments
		STATE_NEXT  = STATE;
		PAUSE_TIME_NEXT = PAUSE_TIME;
		X_PAGE_NEXT = X_PAGE;
		Y_NEXT = Y;
		INDEX_NEXT = INDEX;
		LCD_DI_NEXT = LCD_DI;
		LCD_RW_NEXT = LCD_RW;
		LCD_DATA_NEXT = LCD_DATA;	
		IMAGE_NEXT = IMAGE;
		COL_COUNTER_NEXT = COL_COUNTER; 
		PAGE_COUNTER_NEXT = PAGE_COUNTER;
		START_NEXT =	1'b0;	
		NEW_PAGE_NEXT = 1'b0;
		NEW_COL_NEXT = 1'b0;	
		ENABLE_NEXT = 1'b0;
		//added
		LCD_CS1_NEXT = LCD_CS1;
		LCD_CS2_NEXT = LCD_CS2;
		LCD_SELECT_NEXT = LCD_SELECT;
		LCD_SIDE_NEXT = LCD_SIDE;
		//added
		case(STATE)
			Init: begin  //initial state
				STATE_NEXT =  Set_StartLine;
				// prepare LCD instruction to turn display on
				LCD_DI_NEXT = 1'b0;
				LCD_RW_NEXT = 1'b0;
				LCD_DATA_NEXT = 8'b0011111_1;
				ENABLE_NEXT = 1'b1;
			end
			Set_StartLine: begin //set start line
				STATE_NEXT = Clear_Screen;
				// prepare LCD instruction to set start line
				LCD_DI_NEXT = 1'b0;
				LCD_RW_NEXT = 1'b0;
				LCD_DATA_NEXT = 8'b11_000000; // start line = 0
				ENABLE_NEXT = 1'b1;
				START_NEXT = 1'b1;
			end
			Clear_Screen: begin
				if (START) begin
					NEW_PAGE_NEXT = 1'b1;
					PAGE_COUNTER_NEXT = 0;
					COL_COUNTER_NEXT = 0;
					X_PAGE_NEXT = 0; // set initial X address
					Y_NEXT = 0; // set initial Y address
				end else	
				if (NEW_PAGE) begin
					// prepare LCD instruction to move to new page
					LCD_DI_NEXT = 1'b0;
					LCD_RW_NEXT = 1'd0;
					LCD_DATA_NEXT = {5'b10111, X_PAGE};
					ENABLE_NEXT = 1'b1;
					NEW_COL_NEXT = 1'b1;
				end else if (NEW_COL) begin 
					// prepare LCD instruction to move to column 0 
					LCD_DI_NEXT    = 1'b0;
					LCD_RW_NEXT    = 1'd0;
					LCD_DATA_NEXT  = 8'b01_000000; // to move to column 0
					ENABLE_NEXT = 1'b1;
				end else if (COL_COUNTER < 64) begin
					// prepare LCD instruction to write 00000000 into display RAM
					LCD_DI_NEXT    = 1'b1;
					LCD_RW_NEXT    = 1'd0;
					LCD_DATA_NEXT  = 8'b00000000;
					ENABLE_NEXT = 1'b1;
					COL_COUNTER_NEXT = COL_COUNTER + 1;
				end else begin
					if (PAGE_COUNTER == 7) begin // last page of screen
						STATE_NEXT = Copy_Image;
						START_NEXT = 1'b1;
					end else begin
						// prepare to change page
						X_PAGE_NEXT  = X_PAGE + 1;
						NEW_PAGE_NEXT = 1'b1;
						PAGE_COUNTER_NEXT = PAGE_COUNTER + 1;
						COL_COUNTER_NEXT = 0;
					end
				end
			end						
			Copy_Image: begin // write image pattern into LCD RAM
				if (START) begin
					NEW_PAGE_NEXT = 1'b1;
					X_PAGE_NEXT = 3'b0;  // image initial X address
					Y_NEXT = 0; // image initial Y address
					PAGE_COUNTER_NEXT = 0;
					COL_COUNTER_NEXT = 0;
					//added
					LCD_CS1_NEXT = ~LCD_SELECT;
					LCD_CS2_NEXT = LCD_SELECT;
					//added
				end else if (NEW_PAGE) begin
					// prepare LCD instruction to move to new page 
					LCD_DI_NEXT = 1'b0;
					LCD_RW_NEXT = 1'b0;
					LCD_DATA_NEXT = {5'b10111, X_PAGE}; 
					ENABLE_NEXT = 1'b1;
					NEW_COL_NEXT = 1'b1;
				end else if (NEW_COL) begin
					// prepare LCD instruction to move to new column
					LCD_DI_NEXT = 1'b0;
					LCD_RW_NEXT = 1'b0;
					LCD_DATA_NEXT = {2'b01,Y};
					ENABLE_NEXT = 1'b1;
				end else if (COL_COUNTER < 64) begin //load image 1 byte at a time, 16 is the width of image
					// prepare LCD instruction to write image data into display RAM
					LCD_DI_NEXT = 1'b1;
					LCD_RW_NEXT = 1'b0;
					LCD_DATA_NEXT = PATTERN;
					ENABLE_NEXT = 1'b1;
					INDEX_NEXT = INDEX + 1;
					COL_COUNTER_NEXT = COL_COUNTER + 1;
				end else begin 
					if (PAGE_COUNTER == 7) begin // last page of image
						LCD_SIDE_NEXT = LCD_SIDE + 1;
						if(LCD_SELECT == 0)begin
							LCD_SELECT_NEXT = LCD_SELECT + 1;
							START_NEXT = 1'b1;
						end else if(LCD_SELECT == 1)begin
							LCD_SELECT_NEXT = LCD_SELECT + 1;
							INDEX_NEXT = 0;
							STATE_NEXT = Pause;
						end						
					end else begin
						// prepare to change page
						X_PAGE_NEXT = X_PAGE + 1;		
						NEW_PAGE_NEXT = 1'b1;
						PAGE_COUNTER_NEXT = PAGE_COUNTER + 1;
						COL_COUNTER_NEXT = 0;
					end
				end				
			end
			Pause: begin
				if (PAUSED_TO_THE_END) begin
					STATE_NEXT = Copy_Image;
					START_NEXT = 1'b1;
				end 
				else STATE_NEXT = Pause;
				PAUSE_TIME_NEXT = PAUSE_TIME - 1; 
			end
			default: STATE_NEXT = Init;
		endcase
    end
/******************************
 * Set image patterns		   *
 ******************************/
    always @(*)begin
	case(IMAGE)
		2'b00:	// 1st image 	
			case(LCD_CS1)
				1'b0:
				case (INDEX) // 
				//------PAGE 0-------//
				  	9'd  0	:	PATTERN = {RIGHT_GRAPH[ 448], RIGHT_GRAPH[ 384], RIGHT_GRAPH[ 320], RIGHT_GRAPH[ 256], RIGHT_GRAPH[ 192], RIGHT_GRAPH[ 128], RIGHT_GRAPH[  64], RIGHT_GRAPH[   0]};
					9'd  1	:	PATTERN = {RIGHT_GRAPH[ 449], RIGHT_GRAPH[ 385], RIGHT_GRAPH[ 321], RIGHT_GRAPH[ 257], RIGHT_GRAPH[ 193], RIGHT_GRAPH[ 129], RIGHT_GRAPH[  65], RIGHT_GRAPH[   1]};
					9'd  2	:	PATTERN = {RIGHT_GRAPH[ 450], RIGHT_GRAPH[ 386], RIGHT_GRAPH[ 322], RIGHT_GRAPH[ 258], RIGHT_GRAPH[ 194], RIGHT_GRAPH[ 130], RIGHT_GRAPH[  66], RIGHT_GRAPH[   2]};
					9'd  3	:	PATTERN = {RIGHT_GRAPH[ 451], RIGHT_GRAPH[ 387], RIGHT_GRAPH[ 323], RIGHT_GRAPH[ 259], RIGHT_GRAPH[ 195], RIGHT_GRAPH[ 131], RIGHT_GRAPH[  67], RIGHT_GRAPH[   3]};
					9'd  4	:	PATTERN = {RIGHT_GRAPH[ 452], RIGHT_GRAPH[ 388], RIGHT_GRAPH[ 324], RIGHT_GRAPH[ 260], RIGHT_GRAPH[ 196], RIGHT_GRAPH[ 132], RIGHT_GRAPH[  68], RIGHT_GRAPH[   4]};
					9'd  5	:	PATTERN = {RIGHT_GRAPH[ 453], RIGHT_GRAPH[ 389], RIGHT_GRAPH[ 325], RIGHT_GRAPH[ 261], RIGHT_GRAPH[ 197], RIGHT_GRAPH[ 133], RIGHT_GRAPH[  69], RIGHT_GRAPH[   5]};
					9'd  6	:	PATTERN = {RIGHT_GRAPH[ 454], RIGHT_GRAPH[ 390], RIGHT_GRAPH[ 326], RIGHT_GRAPH[ 262], RIGHT_GRAPH[ 198], RIGHT_GRAPH[ 134], RIGHT_GRAPH[  70], RIGHT_GRAPH[   6]};
					9'd  7	:	PATTERN = {RIGHT_GRAPH[ 455], RIGHT_GRAPH[ 391], RIGHT_GRAPH[ 327], RIGHT_GRAPH[ 263], RIGHT_GRAPH[ 199], RIGHT_GRAPH[ 135], RIGHT_GRAPH[  71], RIGHT_GRAPH[   7]};
					9'd  8	:	PATTERN = {RIGHT_GRAPH[ 456], RIGHT_GRAPH[ 392], RIGHT_GRAPH[ 328], RIGHT_GRAPH[ 264], RIGHT_GRAPH[ 200], RIGHT_GRAPH[ 136], RIGHT_GRAPH[  72], RIGHT_GRAPH[   8]};
					9'd  9	:	PATTERN = {RIGHT_GRAPH[ 457], RIGHT_GRAPH[ 393], RIGHT_GRAPH[ 329], RIGHT_GRAPH[ 265], RIGHT_GRAPH[ 201], RIGHT_GRAPH[ 137], RIGHT_GRAPH[  73], RIGHT_GRAPH[   9]};
					9'd 10	:	PATTERN = {RIGHT_GRAPH[ 458], RIGHT_GRAPH[ 394], RIGHT_GRAPH[ 330], RIGHT_GRAPH[ 266], RIGHT_GRAPH[ 202], RIGHT_GRAPH[ 138], RIGHT_GRAPH[  74], RIGHT_GRAPH[  10]};
					9'd 11	:	PATTERN = {RIGHT_GRAPH[ 459], RIGHT_GRAPH[ 395], RIGHT_GRAPH[ 331], RIGHT_GRAPH[ 267], RIGHT_GRAPH[ 203], RIGHT_GRAPH[ 139], RIGHT_GRAPH[  75], RIGHT_GRAPH[  11]};
					9'd 12	:	PATTERN = {RIGHT_GRAPH[ 460], RIGHT_GRAPH[ 396], RIGHT_GRAPH[ 332], RIGHT_GRAPH[ 268], RIGHT_GRAPH[ 204], RIGHT_GRAPH[ 140], RIGHT_GRAPH[  76], RIGHT_GRAPH[  12]};
					9'd 13	:	PATTERN = {RIGHT_GRAPH[ 461], RIGHT_GRAPH[ 397], RIGHT_GRAPH[ 333], RIGHT_GRAPH[ 269], RIGHT_GRAPH[ 205], RIGHT_GRAPH[ 141], RIGHT_GRAPH[  77], RIGHT_GRAPH[  13]};
					9'd 14	:	PATTERN = {RIGHT_GRAPH[ 462], RIGHT_GRAPH[ 398], RIGHT_GRAPH[ 334], RIGHT_GRAPH[ 270], RIGHT_GRAPH[ 206], RIGHT_GRAPH[ 142], RIGHT_GRAPH[  78], RIGHT_GRAPH[  14]};
					9'd 15	:	PATTERN = {RIGHT_GRAPH[ 463], RIGHT_GRAPH[ 399], RIGHT_GRAPH[ 335], RIGHT_GRAPH[ 271], RIGHT_GRAPH[ 207], RIGHT_GRAPH[ 143], RIGHT_GRAPH[  79], RIGHT_GRAPH[  15]};
					9'd 16	:	PATTERN = {RIGHT_GRAPH[ 464], RIGHT_GRAPH[ 400], RIGHT_GRAPH[ 336], RIGHT_GRAPH[ 272], RIGHT_GRAPH[ 208], RIGHT_GRAPH[ 144], RIGHT_GRAPH[  80], RIGHT_GRAPH[  16]};
					9'd 17	:	PATTERN = {RIGHT_GRAPH[ 465], RIGHT_GRAPH[ 401], RIGHT_GRAPH[ 337], RIGHT_GRAPH[ 273], RIGHT_GRAPH[ 209], RIGHT_GRAPH[ 145], RIGHT_GRAPH[  81], RIGHT_GRAPH[  17]};
					9'd 18	:	PATTERN = {RIGHT_GRAPH[ 466], RIGHT_GRAPH[ 402], RIGHT_GRAPH[ 338], RIGHT_GRAPH[ 274], RIGHT_GRAPH[ 210], RIGHT_GRAPH[ 146], RIGHT_GRAPH[  82], RIGHT_GRAPH[  18]};
					9'd 19	:	PATTERN = {RIGHT_GRAPH[ 467], RIGHT_GRAPH[ 403], RIGHT_GRAPH[ 339], RIGHT_GRAPH[ 275], RIGHT_GRAPH[ 211], RIGHT_GRAPH[ 147], RIGHT_GRAPH[  83], RIGHT_GRAPH[  19]};
					9'd 20	:	PATTERN = {RIGHT_GRAPH[ 468], RIGHT_GRAPH[ 404], RIGHT_GRAPH[ 340], RIGHT_GRAPH[ 276], RIGHT_GRAPH[ 212], RIGHT_GRAPH[ 148], RIGHT_GRAPH[  84], RIGHT_GRAPH[  20]};
					9'd 21	:	PATTERN = {RIGHT_GRAPH[ 469], RIGHT_GRAPH[ 405], RIGHT_GRAPH[ 341], RIGHT_GRAPH[ 277], RIGHT_GRAPH[ 213], RIGHT_GRAPH[ 149], RIGHT_GRAPH[  85], RIGHT_GRAPH[  21]};
					9'd 22	:	PATTERN = {RIGHT_GRAPH[ 470], RIGHT_GRAPH[ 406], RIGHT_GRAPH[ 342], RIGHT_GRAPH[ 278], RIGHT_GRAPH[ 214], RIGHT_GRAPH[ 150], RIGHT_GRAPH[  86], RIGHT_GRAPH[  22]};
					9'd 23	:	PATTERN = {RIGHT_GRAPH[ 471], RIGHT_GRAPH[ 407], RIGHT_GRAPH[ 343], RIGHT_GRAPH[ 279], RIGHT_GRAPH[ 215], RIGHT_GRAPH[ 151], RIGHT_GRAPH[  87], RIGHT_GRAPH[  23]};
					9'd 24	:	PATTERN = {RIGHT_GRAPH[ 472], RIGHT_GRAPH[ 408], RIGHT_GRAPH[ 344], RIGHT_GRAPH[ 280], RIGHT_GRAPH[ 216], RIGHT_GRAPH[ 152], RIGHT_GRAPH[  88], RIGHT_GRAPH[  24]};
					9'd 25	:	PATTERN = {RIGHT_GRAPH[ 473], RIGHT_GRAPH[ 409], RIGHT_GRAPH[ 345], RIGHT_GRAPH[ 281], RIGHT_GRAPH[ 217], RIGHT_GRAPH[ 153], RIGHT_GRAPH[  89], RIGHT_GRAPH[  25]};
					9'd 26	:	PATTERN = {RIGHT_GRAPH[ 474], RIGHT_GRAPH[ 410], RIGHT_GRAPH[ 346], RIGHT_GRAPH[ 282], RIGHT_GRAPH[ 218], RIGHT_GRAPH[ 154], RIGHT_GRAPH[  90], RIGHT_GRAPH[  26]};
					9'd 27	:	PATTERN = {RIGHT_GRAPH[ 475], RIGHT_GRAPH[ 411], RIGHT_GRAPH[ 347], RIGHT_GRAPH[ 283], RIGHT_GRAPH[ 219], RIGHT_GRAPH[ 155], RIGHT_GRAPH[  91], RIGHT_GRAPH[  27]};
					9'd 28	:	PATTERN = {RIGHT_GRAPH[ 476], RIGHT_GRAPH[ 412], RIGHT_GRAPH[ 348], RIGHT_GRAPH[ 284], RIGHT_GRAPH[ 220], RIGHT_GRAPH[ 156], RIGHT_GRAPH[  92], RIGHT_GRAPH[  28]};
					9'd 29	:	PATTERN = {RIGHT_GRAPH[ 477], RIGHT_GRAPH[ 413], RIGHT_GRAPH[ 349], RIGHT_GRAPH[ 285], RIGHT_GRAPH[ 221], RIGHT_GRAPH[ 157], RIGHT_GRAPH[  93], RIGHT_GRAPH[  29]};
					9'd 30	:	PATTERN = {RIGHT_GRAPH[ 478], RIGHT_GRAPH[ 414], RIGHT_GRAPH[ 350], RIGHT_GRAPH[ 286], RIGHT_GRAPH[ 222], RIGHT_GRAPH[ 158], RIGHT_GRAPH[  94], RIGHT_GRAPH[  30]};
					9'd 31	:	PATTERN = {RIGHT_GRAPH[ 479], RIGHT_GRAPH[ 415], RIGHT_GRAPH[ 351], RIGHT_GRAPH[ 287], RIGHT_GRAPH[ 223], RIGHT_GRAPH[ 159], RIGHT_GRAPH[  95], RIGHT_GRAPH[  31]};
					9'd 32	:	PATTERN = {RIGHT_GRAPH[ 480], RIGHT_GRAPH[ 416], RIGHT_GRAPH[ 352], RIGHT_GRAPH[ 288], RIGHT_GRAPH[ 224], RIGHT_GRAPH[ 160], RIGHT_GRAPH[  96], RIGHT_GRAPH[  32]};
					9'd 33	:	PATTERN = {RIGHT_GRAPH[ 481], RIGHT_GRAPH[ 417], RIGHT_GRAPH[ 353], RIGHT_GRAPH[ 289], RIGHT_GRAPH[ 225], RIGHT_GRAPH[ 161], RIGHT_GRAPH[  97], RIGHT_GRAPH[  33]};
					9'd 34	:	PATTERN = {RIGHT_GRAPH[ 482], RIGHT_GRAPH[ 418], RIGHT_GRAPH[ 354], RIGHT_GRAPH[ 290], RIGHT_GRAPH[ 226], RIGHT_GRAPH[ 162], RIGHT_GRAPH[  98], RIGHT_GRAPH[  34]};
					9'd 35	:	PATTERN = {RIGHT_GRAPH[ 483], RIGHT_GRAPH[ 419], RIGHT_GRAPH[ 355], RIGHT_GRAPH[ 291], RIGHT_GRAPH[ 227], RIGHT_GRAPH[ 163], RIGHT_GRAPH[  99], RIGHT_GRAPH[  35]};
					9'd 36	:	PATTERN = {RIGHT_GRAPH[ 484], RIGHT_GRAPH[ 420], RIGHT_GRAPH[ 356], RIGHT_GRAPH[ 292], RIGHT_GRAPH[ 228], RIGHT_GRAPH[ 164], RIGHT_GRAPH[ 100], RIGHT_GRAPH[  36]};
					9'd 37	:	PATTERN = {RIGHT_GRAPH[ 485], RIGHT_GRAPH[ 421], RIGHT_GRAPH[ 357], RIGHT_GRAPH[ 293], RIGHT_GRAPH[ 229], RIGHT_GRAPH[ 165], RIGHT_GRAPH[ 101], RIGHT_GRAPH[  37]};
					9'd 38	:	PATTERN = {RIGHT_GRAPH[ 486], RIGHT_GRAPH[ 422], RIGHT_GRAPH[ 358], RIGHT_GRAPH[ 294], RIGHT_GRAPH[ 230], RIGHT_GRAPH[ 166], RIGHT_GRAPH[ 102], RIGHT_GRAPH[  38]};
					9'd 39	:	PATTERN = {RIGHT_GRAPH[ 487], RIGHT_GRAPH[ 423], RIGHT_GRAPH[ 359], RIGHT_GRAPH[ 295], RIGHT_GRAPH[ 231], RIGHT_GRAPH[ 167], RIGHT_GRAPH[ 103], RIGHT_GRAPH[  39]};
					9'd 40	:	PATTERN = {RIGHT_GRAPH[ 488], RIGHT_GRAPH[ 424], RIGHT_GRAPH[ 360], RIGHT_GRAPH[ 296], RIGHT_GRAPH[ 232], RIGHT_GRAPH[ 168], RIGHT_GRAPH[ 104], RIGHT_GRAPH[  40]};
					9'd 41	:	PATTERN = {RIGHT_GRAPH[ 489], RIGHT_GRAPH[ 425], RIGHT_GRAPH[ 361], RIGHT_GRAPH[ 297], RIGHT_GRAPH[ 233], RIGHT_GRAPH[ 169], RIGHT_GRAPH[ 105], RIGHT_GRAPH[  41]};
					9'd 42	:	PATTERN = {RIGHT_GRAPH[ 490], RIGHT_GRAPH[ 426], RIGHT_GRAPH[ 362], RIGHT_GRAPH[ 298], RIGHT_GRAPH[ 234], RIGHT_GRAPH[ 170], RIGHT_GRAPH[ 106], RIGHT_GRAPH[  42]};
					9'd 43	:	PATTERN = {RIGHT_GRAPH[ 491], RIGHT_GRAPH[ 427], RIGHT_GRAPH[ 363], RIGHT_GRAPH[ 299], RIGHT_GRAPH[ 235], RIGHT_GRAPH[ 171], RIGHT_GRAPH[ 107], RIGHT_GRAPH[  43]};
					9'd 44	:	PATTERN = {RIGHT_GRAPH[ 492], RIGHT_GRAPH[ 428], RIGHT_GRAPH[ 364], RIGHT_GRAPH[ 300], RIGHT_GRAPH[ 236], RIGHT_GRAPH[ 172], RIGHT_GRAPH[ 108], RIGHT_GRAPH[  44]};
					9'd 45	:	PATTERN = {RIGHT_GRAPH[ 493], RIGHT_GRAPH[ 429], RIGHT_GRAPH[ 365], RIGHT_GRAPH[ 301], RIGHT_GRAPH[ 237], RIGHT_GRAPH[ 173], RIGHT_GRAPH[ 109], RIGHT_GRAPH[  45]};
					9'd 46	:	PATTERN = {RIGHT_GRAPH[ 494], RIGHT_GRAPH[ 430], RIGHT_GRAPH[ 366], RIGHT_GRAPH[ 302], RIGHT_GRAPH[ 238], RIGHT_GRAPH[ 174], RIGHT_GRAPH[ 110], RIGHT_GRAPH[  46]};
					9'd 47	:	PATTERN = {RIGHT_GRAPH[ 495], RIGHT_GRAPH[ 431], RIGHT_GRAPH[ 367], RIGHT_GRAPH[ 303], RIGHT_GRAPH[ 239], RIGHT_GRAPH[ 175], RIGHT_GRAPH[ 111], RIGHT_GRAPH[  47]};
					9'd 48	:	PATTERN = {RIGHT_GRAPH[ 496], RIGHT_GRAPH[ 432], RIGHT_GRAPH[ 368], RIGHT_GRAPH[ 304], RIGHT_GRAPH[ 240], RIGHT_GRAPH[ 176], RIGHT_GRAPH[ 112], RIGHT_GRAPH[  48]};
					9'd 49	:	PATTERN = {RIGHT_GRAPH[ 497], RIGHT_GRAPH[ 433], RIGHT_GRAPH[ 369], RIGHT_GRAPH[ 305], RIGHT_GRAPH[ 241], RIGHT_GRAPH[ 177], RIGHT_GRAPH[ 113], RIGHT_GRAPH[  49]};
					9'd 50	:	PATTERN = {RIGHT_GRAPH[ 498], RIGHT_GRAPH[ 434], RIGHT_GRAPH[ 370], RIGHT_GRAPH[ 306], RIGHT_GRAPH[ 242], RIGHT_GRAPH[ 178], RIGHT_GRAPH[ 114], RIGHT_GRAPH[  50]};
					9'd 51	:	PATTERN = {RIGHT_GRAPH[ 499], RIGHT_GRAPH[ 435], RIGHT_GRAPH[ 371], RIGHT_GRAPH[ 307], RIGHT_GRAPH[ 243], RIGHT_GRAPH[ 179], RIGHT_GRAPH[ 115], RIGHT_GRAPH[  51]};
					9'd 52	:	PATTERN = {RIGHT_GRAPH[ 500], RIGHT_GRAPH[ 436], RIGHT_GRAPH[ 372], RIGHT_GRAPH[ 308], RIGHT_GRAPH[ 244], RIGHT_GRAPH[ 180], RIGHT_GRAPH[ 116], RIGHT_GRAPH[  52]};
					9'd 53	:	PATTERN = {RIGHT_GRAPH[ 501], RIGHT_GRAPH[ 437], RIGHT_GRAPH[ 373], RIGHT_GRAPH[ 309], RIGHT_GRAPH[ 245], RIGHT_GRAPH[ 181], RIGHT_GRAPH[ 117], RIGHT_GRAPH[  53]};
					9'd 54	:	PATTERN = {RIGHT_GRAPH[ 502], RIGHT_GRAPH[ 438], RIGHT_GRAPH[ 374], RIGHT_GRAPH[ 310], RIGHT_GRAPH[ 246], RIGHT_GRAPH[ 182], RIGHT_GRAPH[ 118], RIGHT_GRAPH[  54]};
					9'd 55	:	PATTERN = {RIGHT_GRAPH[ 503], RIGHT_GRAPH[ 439], RIGHT_GRAPH[ 375], RIGHT_GRAPH[ 311], RIGHT_GRAPH[ 247], RIGHT_GRAPH[ 183], RIGHT_GRAPH[ 119], RIGHT_GRAPH[  55]};
					9'd 56	:	PATTERN = {RIGHT_GRAPH[ 504], RIGHT_GRAPH[ 440], RIGHT_GRAPH[ 376], RIGHT_GRAPH[ 312], RIGHT_GRAPH[ 248], RIGHT_GRAPH[ 184], RIGHT_GRAPH[ 120], RIGHT_GRAPH[  56]};
					9'd 57	:	PATTERN = {RIGHT_GRAPH[ 505], RIGHT_GRAPH[ 441], RIGHT_GRAPH[ 377], RIGHT_GRAPH[ 313], RIGHT_GRAPH[ 249], RIGHT_GRAPH[ 185], RIGHT_GRAPH[ 121], RIGHT_GRAPH[  57]};
					9'd 58	:	PATTERN = {RIGHT_GRAPH[ 506], RIGHT_GRAPH[ 442], RIGHT_GRAPH[ 378], RIGHT_GRAPH[ 314], RIGHT_GRAPH[ 250], RIGHT_GRAPH[ 186], RIGHT_GRAPH[ 122], RIGHT_GRAPH[  58]};
					9'd 59	:	PATTERN = {RIGHT_GRAPH[ 507], RIGHT_GRAPH[ 443], RIGHT_GRAPH[ 379], RIGHT_GRAPH[ 315], RIGHT_GRAPH[ 251], RIGHT_GRAPH[ 187], RIGHT_GRAPH[ 123], RIGHT_GRAPH[  59]};
					9'd 60	:	PATTERN = {RIGHT_GRAPH[ 508], RIGHT_GRAPH[ 444], RIGHT_GRAPH[ 380], RIGHT_GRAPH[ 316], RIGHT_GRAPH[ 252], RIGHT_GRAPH[ 188], RIGHT_GRAPH[ 124], RIGHT_GRAPH[  60]};
					9'd 61	:	PATTERN = {RIGHT_GRAPH[ 509], RIGHT_GRAPH[ 445], RIGHT_GRAPH[ 381], RIGHT_GRAPH[ 317], RIGHT_GRAPH[ 253], RIGHT_GRAPH[ 189], RIGHT_GRAPH[ 125], RIGHT_GRAPH[  61]};
					9'd 62	:	PATTERN = {RIGHT_GRAPH[ 510], RIGHT_GRAPH[ 446], RIGHT_GRAPH[ 382], RIGHT_GRAPH[ 318], RIGHT_GRAPH[ 254], RIGHT_GRAPH[ 190], RIGHT_GRAPH[ 126], RIGHT_GRAPH[  62]};
					9'd 63	:	PATTERN = {RIGHT_GRAPH[ 511], RIGHT_GRAPH[ 447], RIGHT_GRAPH[ 383], RIGHT_GRAPH[ 319], RIGHT_GRAPH[ 255], RIGHT_GRAPH[ 191], RIGHT_GRAPH[ 127], RIGHT_GRAPH[  63]};
					9'd 64	:	PATTERN = {RIGHT_GRAPH[ 960], RIGHT_GRAPH[ 896], RIGHT_GRAPH[ 832], RIGHT_GRAPH[ 768], RIGHT_GRAPH[ 704], RIGHT_GRAPH[ 640], RIGHT_GRAPH[ 576], RIGHT_GRAPH[ 512]};
					9'd 65	:	PATTERN = {RIGHT_GRAPH[ 961], RIGHT_GRAPH[ 897], RIGHT_GRAPH[ 833], RIGHT_GRAPH[ 769], RIGHT_GRAPH[ 705], RIGHT_GRAPH[ 641], RIGHT_GRAPH[ 577], RIGHT_GRAPH[ 513]};
					9'd 66	:	PATTERN = {RIGHT_GRAPH[ 962], RIGHT_GRAPH[ 898], RIGHT_GRAPH[ 834], RIGHT_GRAPH[ 770], RIGHT_GRAPH[ 706], RIGHT_GRAPH[ 642], RIGHT_GRAPH[ 578], RIGHT_GRAPH[ 514]};
					9'd 67	:	PATTERN = {RIGHT_GRAPH[ 963], RIGHT_GRAPH[ 899], RIGHT_GRAPH[ 835], RIGHT_GRAPH[ 771], RIGHT_GRAPH[ 707], RIGHT_GRAPH[ 643], RIGHT_GRAPH[ 579], RIGHT_GRAPH[ 515]};
					9'd 68	:	PATTERN = {RIGHT_GRAPH[ 964], RIGHT_GRAPH[ 900], RIGHT_GRAPH[ 836], RIGHT_GRAPH[ 772], RIGHT_GRAPH[ 708], RIGHT_GRAPH[ 644], RIGHT_GRAPH[ 580], RIGHT_GRAPH[ 516]};
					9'd 69	:	PATTERN = {RIGHT_GRAPH[ 965], RIGHT_GRAPH[ 901], RIGHT_GRAPH[ 837], RIGHT_GRAPH[ 773], RIGHT_GRAPH[ 709], RIGHT_GRAPH[ 645], RIGHT_GRAPH[ 581], RIGHT_GRAPH[ 517]};
					9'd 70	:	PATTERN = {RIGHT_GRAPH[ 966], RIGHT_GRAPH[ 902], RIGHT_GRAPH[ 838], RIGHT_GRAPH[ 774], RIGHT_GRAPH[ 710], RIGHT_GRAPH[ 646], RIGHT_GRAPH[ 582], RIGHT_GRAPH[ 518]};
					9'd 71	:	PATTERN = {RIGHT_GRAPH[ 967], RIGHT_GRAPH[ 903], RIGHT_GRAPH[ 839], RIGHT_GRAPH[ 775], RIGHT_GRAPH[ 711], RIGHT_GRAPH[ 647], RIGHT_GRAPH[ 583], RIGHT_GRAPH[ 519]};
					9'd 72	:	PATTERN = {RIGHT_GRAPH[ 968], RIGHT_GRAPH[ 904], RIGHT_GRAPH[ 840], RIGHT_GRAPH[ 776], RIGHT_GRAPH[ 712], RIGHT_GRAPH[ 648], RIGHT_GRAPH[ 584], RIGHT_GRAPH[ 520]};
					9'd 73	:	PATTERN = {RIGHT_GRAPH[ 969], RIGHT_GRAPH[ 905], RIGHT_GRAPH[ 841], RIGHT_GRAPH[ 777], RIGHT_GRAPH[ 713], RIGHT_GRAPH[ 649], RIGHT_GRAPH[ 585], RIGHT_GRAPH[ 521]};
					9'd 74	:	PATTERN = {RIGHT_GRAPH[ 970], RIGHT_GRAPH[ 906], RIGHT_GRAPH[ 842], RIGHT_GRAPH[ 778], RIGHT_GRAPH[ 714], RIGHT_GRAPH[ 650], RIGHT_GRAPH[ 586], RIGHT_GRAPH[ 522]};
					9'd 75	:	PATTERN = {RIGHT_GRAPH[ 971], RIGHT_GRAPH[ 907], RIGHT_GRAPH[ 843], RIGHT_GRAPH[ 779], RIGHT_GRAPH[ 715], RIGHT_GRAPH[ 651], RIGHT_GRAPH[ 587], RIGHT_GRAPH[ 523]};
					9'd 76	:	PATTERN = {RIGHT_GRAPH[ 972], RIGHT_GRAPH[ 908], RIGHT_GRAPH[ 844], RIGHT_GRAPH[ 780], RIGHT_GRAPH[ 716], RIGHT_GRAPH[ 652], RIGHT_GRAPH[ 588], RIGHT_GRAPH[ 524]};
					9'd 77	:	PATTERN = {RIGHT_GRAPH[ 973], RIGHT_GRAPH[ 909], RIGHT_GRAPH[ 845], RIGHT_GRAPH[ 781], RIGHT_GRAPH[ 717], RIGHT_GRAPH[ 653], RIGHT_GRAPH[ 589], RIGHT_GRAPH[ 525]};
					9'd 78	:	PATTERN = {RIGHT_GRAPH[ 974], RIGHT_GRAPH[ 910], RIGHT_GRAPH[ 846], RIGHT_GRAPH[ 782], RIGHT_GRAPH[ 718], RIGHT_GRAPH[ 654], RIGHT_GRAPH[ 590], RIGHT_GRAPH[ 526]};
					9'd 79	:	PATTERN = {RIGHT_GRAPH[ 975], RIGHT_GRAPH[ 911], RIGHT_GRAPH[ 847], RIGHT_GRAPH[ 783], RIGHT_GRAPH[ 719], RIGHT_GRAPH[ 655], RIGHT_GRAPH[ 591], RIGHT_GRAPH[ 527]};
					9'd 80	:	PATTERN = {RIGHT_GRAPH[ 976], RIGHT_GRAPH[ 912], RIGHT_GRAPH[ 848], RIGHT_GRAPH[ 784], RIGHT_GRAPH[ 720], RIGHT_GRAPH[ 656], RIGHT_GRAPH[ 592], RIGHT_GRAPH[ 528]};
					9'd 81	:	PATTERN = {RIGHT_GRAPH[ 977], RIGHT_GRAPH[ 913], RIGHT_GRAPH[ 849], RIGHT_GRAPH[ 785], RIGHT_GRAPH[ 721], RIGHT_GRAPH[ 657], RIGHT_GRAPH[ 593], RIGHT_GRAPH[ 529]};
					9'd 82	:	PATTERN = {RIGHT_GRAPH[ 978], RIGHT_GRAPH[ 914], RIGHT_GRAPH[ 850], RIGHT_GRAPH[ 786], RIGHT_GRAPH[ 722], RIGHT_GRAPH[ 658], RIGHT_GRAPH[ 594], RIGHT_GRAPH[ 530]};
					9'd 83	:	PATTERN = {RIGHT_GRAPH[ 979], RIGHT_GRAPH[ 915], RIGHT_GRAPH[ 851], RIGHT_GRAPH[ 787], RIGHT_GRAPH[ 723], RIGHT_GRAPH[ 659], RIGHT_GRAPH[ 595], RIGHT_GRAPH[ 531]};
					9'd 84	:	PATTERN = {RIGHT_GRAPH[ 980], RIGHT_GRAPH[ 916], RIGHT_GRAPH[ 852], RIGHT_GRAPH[ 788], RIGHT_GRAPH[ 724], RIGHT_GRAPH[ 660], RIGHT_GRAPH[ 596], RIGHT_GRAPH[ 532]};
					9'd 85	:	PATTERN = {RIGHT_GRAPH[ 981], RIGHT_GRAPH[ 917], RIGHT_GRAPH[ 853], RIGHT_GRAPH[ 789], RIGHT_GRAPH[ 725], RIGHT_GRAPH[ 661], RIGHT_GRAPH[ 597], RIGHT_GRAPH[ 533]};
					9'd 86	:	PATTERN = {RIGHT_GRAPH[ 982], RIGHT_GRAPH[ 918], RIGHT_GRAPH[ 854], RIGHT_GRAPH[ 790], RIGHT_GRAPH[ 726], RIGHT_GRAPH[ 662], RIGHT_GRAPH[ 598], RIGHT_GRAPH[ 534]};
					9'd 87	:	PATTERN = {RIGHT_GRAPH[ 983], RIGHT_GRAPH[ 919], RIGHT_GRAPH[ 855], RIGHT_GRAPH[ 791], RIGHT_GRAPH[ 727], RIGHT_GRAPH[ 663], RIGHT_GRAPH[ 599], RIGHT_GRAPH[ 535]};
					9'd 88	:	PATTERN = {RIGHT_GRAPH[ 984], RIGHT_GRAPH[ 920], RIGHT_GRAPH[ 856], RIGHT_GRAPH[ 792], RIGHT_GRAPH[ 728], RIGHT_GRAPH[ 664], RIGHT_GRAPH[ 600], RIGHT_GRAPH[ 536]};
					9'd 89	:	PATTERN = {RIGHT_GRAPH[ 985], RIGHT_GRAPH[ 921], RIGHT_GRAPH[ 857], RIGHT_GRAPH[ 793], RIGHT_GRAPH[ 729], RIGHT_GRAPH[ 665], RIGHT_GRAPH[ 601], RIGHT_GRAPH[ 537]};
					9'd 90	:	PATTERN = {RIGHT_GRAPH[ 986], RIGHT_GRAPH[ 922], RIGHT_GRAPH[ 858], RIGHT_GRAPH[ 794], RIGHT_GRAPH[ 730], RIGHT_GRAPH[ 666], RIGHT_GRAPH[ 602], RIGHT_GRAPH[ 538]};
					9'd 91	:	PATTERN = {RIGHT_GRAPH[ 987], RIGHT_GRAPH[ 923], RIGHT_GRAPH[ 859], RIGHT_GRAPH[ 795], RIGHT_GRAPH[ 731], RIGHT_GRAPH[ 667], RIGHT_GRAPH[ 603], RIGHT_GRAPH[ 539]};
					9'd 92	:	PATTERN = {RIGHT_GRAPH[ 988], RIGHT_GRAPH[ 924], RIGHT_GRAPH[ 860], RIGHT_GRAPH[ 796], RIGHT_GRAPH[ 732], RIGHT_GRAPH[ 668], RIGHT_GRAPH[ 604], RIGHT_GRAPH[ 540]};
					9'd 93	:	PATTERN = {RIGHT_GRAPH[ 989], RIGHT_GRAPH[ 925], RIGHT_GRAPH[ 861], RIGHT_GRAPH[ 797], RIGHT_GRAPH[ 733], RIGHT_GRAPH[ 669], RIGHT_GRAPH[ 605], RIGHT_GRAPH[ 541]};
					9'd 94	:	PATTERN = {RIGHT_GRAPH[ 990], RIGHT_GRAPH[ 926], RIGHT_GRAPH[ 862], RIGHT_GRAPH[ 798], RIGHT_GRAPH[ 734], RIGHT_GRAPH[ 670], RIGHT_GRAPH[ 606], RIGHT_GRAPH[ 542]};
					9'd 95	:	PATTERN = {RIGHT_GRAPH[ 991], RIGHT_GRAPH[ 927], RIGHT_GRAPH[ 863], RIGHT_GRAPH[ 799], RIGHT_GRAPH[ 735], RIGHT_GRAPH[ 671], RIGHT_GRAPH[ 607], RIGHT_GRAPH[ 543]};
					9'd 96	:	PATTERN = {RIGHT_GRAPH[ 992], RIGHT_GRAPH[ 928], RIGHT_GRAPH[ 864], RIGHT_GRAPH[ 800], RIGHT_GRAPH[ 736], RIGHT_GRAPH[ 672], RIGHT_GRAPH[ 608], RIGHT_GRAPH[ 544]};
					9'd 97	:	PATTERN = {RIGHT_GRAPH[ 993], RIGHT_GRAPH[ 929], RIGHT_GRAPH[ 865], RIGHT_GRAPH[ 801], RIGHT_GRAPH[ 737], RIGHT_GRAPH[ 673], RIGHT_GRAPH[ 609], RIGHT_GRAPH[ 545]};
					9'd 98	:	PATTERN = {RIGHT_GRAPH[ 994], RIGHT_GRAPH[ 930], RIGHT_GRAPH[ 866], RIGHT_GRAPH[ 802], RIGHT_GRAPH[ 738], RIGHT_GRAPH[ 674], RIGHT_GRAPH[ 610], RIGHT_GRAPH[ 546]};
					9'd 99	:	PATTERN = {RIGHT_GRAPH[ 995], RIGHT_GRAPH[ 931], RIGHT_GRAPH[ 867], RIGHT_GRAPH[ 803], RIGHT_GRAPH[ 739], RIGHT_GRAPH[ 675], RIGHT_GRAPH[ 611], RIGHT_GRAPH[ 547]};
					9'd100	:	PATTERN = {RIGHT_GRAPH[ 996], RIGHT_GRAPH[ 932], RIGHT_GRAPH[ 868], RIGHT_GRAPH[ 804], RIGHT_GRAPH[ 740], RIGHT_GRAPH[ 676], RIGHT_GRAPH[ 612], RIGHT_GRAPH[ 548]};
					9'd101	:	PATTERN = {RIGHT_GRAPH[ 997], RIGHT_GRAPH[ 933], RIGHT_GRAPH[ 869], RIGHT_GRAPH[ 805], RIGHT_GRAPH[ 741], RIGHT_GRAPH[ 677], RIGHT_GRAPH[ 613], RIGHT_GRAPH[ 549]};
					9'd102	:	PATTERN = {RIGHT_GRAPH[ 998], RIGHT_GRAPH[ 934], RIGHT_GRAPH[ 870], RIGHT_GRAPH[ 806], RIGHT_GRAPH[ 742], RIGHT_GRAPH[ 678], RIGHT_GRAPH[ 614], RIGHT_GRAPH[ 550]};
					9'd103	:	PATTERN = {RIGHT_GRAPH[ 999], RIGHT_GRAPH[ 935], RIGHT_GRAPH[ 871], RIGHT_GRAPH[ 807], RIGHT_GRAPH[ 743], RIGHT_GRAPH[ 679], RIGHT_GRAPH[ 615], RIGHT_GRAPH[ 551]};
					9'd104	:	PATTERN = {RIGHT_GRAPH[1000], RIGHT_GRAPH[ 936], RIGHT_GRAPH[ 872], RIGHT_GRAPH[ 808], RIGHT_GRAPH[ 744], RIGHT_GRAPH[ 680], RIGHT_GRAPH[ 616], RIGHT_GRAPH[ 552]};
					9'd105	:	PATTERN = {RIGHT_GRAPH[1001], RIGHT_GRAPH[ 937], RIGHT_GRAPH[ 873], RIGHT_GRAPH[ 809], RIGHT_GRAPH[ 745], RIGHT_GRAPH[ 681], RIGHT_GRAPH[ 617], RIGHT_GRAPH[ 553]};
					9'd106	:	PATTERN = {RIGHT_GRAPH[1002], RIGHT_GRAPH[ 938], RIGHT_GRAPH[ 874], RIGHT_GRAPH[ 810], RIGHT_GRAPH[ 746], RIGHT_GRAPH[ 682], RIGHT_GRAPH[ 618], RIGHT_GRAPH[ 554]};
					9'd107	:	PATTERN = {RIGHT_GRAPH[1003], RIGHT_GRAPH[ 939], RIGHT_GRAPH[ 875], RIGHT_GRAPH[ 811], RIGHT_GRAPH[ 747], RIGHT_GRAPH[ 683], RIGHT_GRAPH[ 619], RIGHT_GRAPH[ 555]};
					9'd108	:	PATTERN = {RIGHT_GRAPH[1004], RIGHT_GRAPH[ 940], RIGHT_GRAPH[ 876], RIGHT_GRAPH[ 812], RIGHT_GRAPH[ 748], RIGHT_GRAPH[ 684], RIGHT_GRAPH[ 620], RIGHT_GRAPH[ 556]};
					9'd109	:	PATTERN = {RIGHT_GRAPH[1005], RIGHT_GRAPH[ 941], RIGHT_GRAPH[ 877], RIGHT_GRAPH[ 813], RIGHT_GRAPH[ 749], RIGHT_GRAPH[ 685], RIGHT_GRAPH[ 621], RIGHT_GRAPH[ 557]};
					9'd110	:	PATTERN = {RIGHT_GRAPH[1006], RIGHT_GRAPH[ 942], RIGHT_GRAPH[ 878], RIGHT_GRAPH[ 814], RIGHT_GRAPH[ 750], RIGHT_GRAPH[ 686], RIGHT_GRAPH[ 622], RIGHT_GRAPH[ 558]};
					9'd111	:	PATTERN = {RIGHT_GRAPH[1007], RIGHT_GRAPH[ 943], RIGHT_GRAPH[ 879], RIGHT_GRAPH[ 815], RIGHT_GRAPH[ 751], RIGHT_GRAPH[ 687], RIGHT_GRAPH[ 623], RIGHT_GRAPH[ 559]};
					9'd112	:	PATTERN = {RIGHT_GRAPH[1008], RIGHT_GRAPH[ 944], RIGHT_GRAPH[ 880], RIGHT_GRAPH[ 816], RIGHT_GRAPH[ 752], RIGHT_GRAPH[ 688], RIGHT_GRAPH[ 624], RIGHT_GRAPH[ 560]};
					9'd113	:	PATTERN = {RIGHT_GRAPH[1009], RIGHT_GRAPH[ 945], RIGHT_GRAPH[ 881], RIGHT_GRAPH[ 817], RIGHT_GRAPH[ 753], RIGHT_GRAPH[ 689], RIGHT_GRAPH[ 625], RIGHT_GRAPH[ 561]};
					9'd114	:	PATTERN = {RIGHT_GRAPH[1010], RIGHT_GRAPH[ 946], RIGHT_GRAPH[ 882], RIGHT_GRAPH[ 818], RIGHT_GRAPH[ 754], RIGHT_GRAPH[ 690], RIGHT_GRAPH[ 626], RIGHT_GRAPH[ 562]};
					9'd115	:	PATTERN = {RIGHT_GRAPH[1011], RIGHT_GRAPH[ 947], RIGHT_GRAPH[ 883], RIGHT_GRAPH[ 819], RIGHT_GRAPH[ 755], RIGHT_GRAPH[ 691], RIGHT_GRAPH[ 627], RIGHT_GRAPH[ 563]};
					9'd116	:	PATTERN = {RIGHT_GRAPH[1012], RIGHT_GRAPH[ 948], RIGHT_GRAPH[ 884], RIGHT_GRAPH[ 820], RIGHT_GRAPH[ 756], RIGHT_GRAPH[ 692], RIGHT_GRAPH[ 628], RIGHT_GRAPH[ 564]};
					9'd117	:	PATTERN = {RIGHT_GRAPH[1013], RIGHT_GRAPH[ 949], RIGHT_GRAPH[ 885], RIGHT_GRAPH[ 821], RIGHT_GRAPH[ 757], RIGHT_GRAPH[ 693], RIGHT_GRAPH[ 629], RIGHT_GRAPH[ 565]};
					9'd118	:	PATTERN = {RIGHT_GRAPH[1014], RIGHT_GRAPH[ 950], RIGHT_GRAPH[ 886], RIGHT_GRAPH[ 822], RIGHT_GRAPH[ 758], RIGHT_GRAPH[ 694], RIGHT_GRAPH[ 630], RIGHT_GRAPH[ 566]};
					9'd119	:	PATTERN = {RIGHT_GRAPH[1015], RIGHT_GRAPH[ 951], RIGHT_GRAPH[ 887], RIGHT_GRAPH[ 823], RIGHT_GRAPH[ 759], RIGHT_GRAPH[ 695], RIGHT_GRAPH[ 631], RIGHT_GRAPH[ 567]};
					9'd120	:	PATTERN = {RIGHT_GRAPH[1016], RIGHT_GRAPH[ 952], RIGHT_GRAPH[ 888], RIGHT_GRAPH[ 824], RIGHT_GRAPH[ 760], RIGHT_GRAPH[ 696], RIGHT_GRAPH[ 632], RIGHT_GRAPH[ 568]};
					9'd121	:	PATTERN = {RIGHT_GRAPH[1017], RIGHT_GRAPH[ 953], RIGHT_GRAPH[ 889], RIGHT_GRAPH[ 825], RIGHT_GRAPH[ 761], RIGHT_GRAPH[ 697], RIGHT_GRAPH[ 633], RIGHT_GRAPH[ 569]};
					9'd122	:	PATTERN = {RIGHT_GRAPH[1018], RIGHT_GRAPH[ 954], RIGHT_GRAPH[ 890], RIGHT_GRAPH[ 826], RIGHT_GRAPH[ 762], RIGHT_GRAPH[ 698], RIGHT_GRAPH[ 634], RIGHT_GRAPH[ 570]};
					9'd123	:	PATTERN = {RIGHT_GRAPH[1019], RIGHT_GRAPH[ 955], RIGHT_GRAPH[ 891], RIGHT_GRAPH[ 827], RIGHT_GRAPH[ 763], RIGHT_GRAPH[ 699], RIGHT_GRAPH[ 635], RIGHT_GRAPH[ 571]};
					9'd124	:	PATTERN = {RIGHT_GRAPH[1020], RIGHT_GRAPH[ 956], RIGHT_GRAPH[ 892], RIGHT_GRAPH[ 828], RIGHT_GRAPH[ 764], RIGHT_GRAPH[ 700], RIGHT_GRAPH[ 636], RIGHT_GRAPH[ 572]};
					9'd125	:	PATTERN = {RIGHT_GRAPH[1021], RIGHT_GRAPH[ 957], RIGHT_GRAPH[ 893], RIGHT_GRAPH[ 829], RIGHT_GRAPH[ 765], RIGHT_GRAPH[ 701], RIGHT_GRAPH[ 637], RIGHT_GRAPH[ 573]};
					9'd126	:	PATTERN = {RIGHT_GRAPH[1022], RIGHT_GRAPH[ 958], RIGHT_GRAPH[ 894], RIGHT_GRAPH[ 830], RIGHT_GRAPH[ 766], RIGHT_GRAPH[ 702], RIGHT_GRAPH[ 638], RIGHT_GRAPH[ 574]};
					9'd127	:	PATTERN = {RIGHT_GRAPH[1023], RIGHT_GRAPH[ 959], RIGHT_GRAPH[ 895], RIGHT_GRAPH[ 831], RIGHT_GRAPH[ 767], RIGHT_GRAPH[ 703], RIGHT_GRAPH[ 639], RIGHT_GRAPH[ 575]};
					9'd128	:	PATTERN = {RIGHT_GRAPH[1472], RIGHT_GRAPH[1408], RIGHT_GRAPH[1344], RIGHT_GRAPH[1280], RIGHT_GRAPH[1216], RIGHT_GRAPH[1152], RIGHT_GRAPH[1088], RIGHT_GRAPH[1024]};
					9'd129	:	PATTERN = {RIGHT_GRAPH[1473], RIGHT_GRAPH[1409], RIGHT_GRAPH[1345], RIGHT_GRAPH[1281], RIGHT_GRAPH[1217], RIGHT_GRAPH[1153], RIGHT_GRAPH[1089], RIGHT_GRAPH[1025]};
					9'd130	:	PATTERN = {RIGHT_GRAPH[1474], RIGHT_GRAPH[1410], RIGHT_GRAPH[1346], RIGHT_GRAPH[1282], RIGHT_GRAPH[1218], RIGHT_GRAPH[1154], RIGHT_GRAPH[1090], RIGHT_GRAPH[1026]};
					9'd131	:	PATTERN = {RIGHT_GRAPH[1475], RIGHT_GRAPH[1411], RIGHT_GRAPH[1347], RIGHT_GRAPH[1283], RIGHT_GRAPH[1219], RIGHT_GRAPH[1155], RIGHT_GRAPH[1091], RIGHT_GRAPH[1027]};
					9'd132	:	PATTERN = {RIGHT_GRAPH[1476], RIGHT_GRAPH[1412], RIGHT_GRAPH[1348], RIGHT_GRAPH[1284], RIGHT_GRAPH[1220], RIGHT_GRAPH[1156], RIGHT_GRAPH[1092], RIGHT_GRAPH[1028]};
					9'd133	:	PATTERN = {RIGHT_GRAPH[1477], RIGHT_GRAPH[1413], RIGHT_GRAPH[1349], RIGHT_GRAPH[1285], RIGHT_GRAPH[1221], RIGHT_GRAPH[1157], RIGHT_GRAPH[1093], RIGHT_GRAPH[1029]};
					9'd134	:	PATTERN = {RIGHT_GRAPH[1478], RIGHT_GRAPH[1414], RIGHT_GRAPH[1350], RIGHT_GRAPH[1286], RIGHT_GRAPH[1222], RIGHT_GRAPH[1158], RIGHT_GRAPH[1094], RIGHT_GRAPH[1030]};
					9'd135	:	PATTERN = {RIGHT_GRAPH[1479], RIGHT_GRAPH[1415], RIGHT_GRAPH[1351], RIGHT_GRAPH[1287], RIGHT_GRAPH[1223], RIGHT_GRAPH[1159], RIGHT_GRAPH[1095], RIGHT_GRAPH[1031]};
					9'd136	:	PATTERN = {RIGHT_GRAPH[1480], RIGHT_GRAPH[1416], RIGHT_GRAPH[1352], RIGHT_GRAPH[1288], RIGHT_GRAPH[1224], RIGHT_GRAPH[1160], RIGHT_GRAPH[1096], RIGHT_GRAPH[1032]};
					9'd137	:	PATTERN = {RIGHT_GRAPH[1481], RIGHT_GRAPH[1417], RIGHT_GRAPH[1353], RIGHT_GRAPH[1289], RIGHT_GRAPH[1225], RIGHT_GRAPH[1161], RIGHT_GRAPH[1097], RIGHT_GRAPH[1033]};
					9'd138	:	PATTERN = {RIGHT_GRAPH[1482], RIGHT_GRAPH[1418], RIGHT_GRAPH[1354], RIGHT_GRAPH[1290], RIGHT_GRAPH[1226], RIGHT_GRAPH[1162], RIGHT_GRAPH[1098], RIGHT_GRAPH[1034]};
					9'd139	:	PATTERN = {RIGHT_GRAPH[1483], RIGHT_GRAPH[1419], RIGHT_GRAPH[1355], RIGHT_GRAPH[1291], RIGHT_GRAPH[1227], RIGHT_GRAPH[1163], RIGHT_GRAPH[1099], RIGHT_GRAPH[1035]};
					9'd140	:	PATTERN = {RIGHT_GRAPH[1484], RIGHT_GRAPH[1420], RIGHT_GRAPH[1356], RIGHT_GRAPH[1292], RIGHT_GRAPH[1228], RIGHT_GRAPH[1164], RIGHT_GRAPH[1100], RIGHT_GRAPH[1036]};
					9'd141	:	PATTERN = {RIGHT_GRAPH[1485], RIGHT_GRAPH[1421], RIGHT_GRAPH[1357], RIGHT_GRAPH[1293], RIGHT_GRAPH[1229], RIGHT_GRAPH[1165], RIGHT_GRAPH[1101], RIGHT_GRAPH[1037]};
					9'd142	:	PATTERN = {RIGHT_GRAPH[1486], RIGHT_GRAPH[1422], RIGHT_GRAPH[1358], RIGHT_GRAPH[1294], RIGHT_GRAPH[1230], RIGHT_GRAPH[1166], RIGHT_GRAPH[1102], RIGHT_GRAPH[1038]};
					9'd143	:	PATTERN = {RIGHT_GRAPH[1487], RIGHT_GRAPH[1423], RIGHT_GRAPH[1359], RIGHT_GRAPH[1295], RIGHT_GRAPH[1231], RIGHT_GRAPH[1167], RIGHT_GRAPH[1103], RIGHT_GRAPH[1039]};
					9'd144	:	PATTERN = {RIGHT_GRAPH[1488], RIGHT_GRAPH[1424], RIGHT_GRAPH[1360], RIGHT_GRAPH[1296], RIGHT_GRAPH[1232], RIGHT_GRAPH[1168], RIGHT_GRAPH[1104], RIGHT_GRAPH[1040]};
					9'd145	:	PATTERN = {RIGHT_GRAPH[1489], RIGHT_GRAPH[1425], RIGHT_GRAPH[1361], RIGHT_GRAPH[1297], RIGHT_GRAPH[1233], RIGHT_GRAPH[1169], RIGHT_GRAPH[1105], RIGHT_GRAPH[1041]};
					9'd146	:	PATTERN = {RIGHT_GRAPH[1490], RIGHT_GRAPH[1426], RIGHT_GRAPH[1362], RIGHT_GRAPH[1298], RIGHT_GRAPH[1234], RIGHT_GRAPH[1170], RIGHT_GRAPH[1106], RIGHT_GRAPH[1042]};
					9'd147	:	PATTERN = {RIGHT_GRAPH[1491], RIGHT_GRAPH[1427], RIGHT_GRAPH[1363], RIGHT_GRAPH[1299], RIGHT_GRAPH[1235], RIGHT_GRAPH[1171], RIGHT_GRAPH[1107], RIGHT_GRAPH[1043]};
					9'd148	:	PATTERN = {RIGHT_GRAPH[1492], RIGHT_GRAPH[1428], RIGHT_GRAPH[1364], RIGHT_GRAPH[1300], RIGHT_GRAPH[1236], RIGHT_GRAPH[1172], RIGHT_GRAPH[1108], RIGHT_GRAPH[1044]};
					9'd149	:	PATTERN = {RIGHT_GRAPH[1493], RIGHT_GRAPH[1429], RIGHT_GRAPH[1365], RIGHT_GRAPH[1301], RIGHT_GRAPH[1237], RIGHT_GRAPH[1173], RIGHT_GRAPH[1109], RIGHT_GRAPH[1045]};
					9'd150	:	PATTERN = {RIGHT_GRAPH[1494], RIGHT_GRAPH[1430], RIGHT_GRAPH[1366], RIGHT_GRAPH[1302], RIGHT_GRAPH[1238], RIGHT_GRAPH[1174], RIGHT_GRAPH[1110], RIGHT_GRAPH[1046]};
					9'd151	:	PATTERN = {RIGHT_GRAPH[1495], RIGHT_GRAPH[1431], RIGHT_GRAPH[1367], RIGHT_GRAPH[1303], RIGHT_GRAPH[1239], RIGHT_GRAPH[1175], RIGHT_GRAPH[1111], RIGHT_GRAPH[1047]};
					9'd152	:	PATTERN = {RIGHT_GRAPH[1496], RIGHT_GRAPH[1432], RIGHT_GRAPH[1368], RIGHT_GRAPH[1304], RIGHT_GRAPH[1240], RIGHT_GRAPH[1176], RIGHT_GRAPH[1112], RIGHT_GRAPH[1048]};
					9'd153	:	PATTERN = {RIGHT_GRAPH[1497], RIGHT_GRAPH[1433], RIGHT_GRAPH[1369], RIGHT_GRAPH[1305], RIGHT_GRAPH[1241], RIGHT_GRAPH[1177], RIGHT_GRAPH[1113], RIGHT_GRAPH[1049]};
					9'd154	:	PATTERN = {RIGHT_GRAPH[1498], RIGHT_GRAPH[1434], RIGHT_GRAPH[1370], RIGHT_GRAPH[1306], RIGHT_GRAPH[1242], RIGHT_GRAPH[1178], RIGHT_GRAPH[1114], RIGHT_GRAPH[1050]};
					9'd155	:	PATTERN = {RIGHT_GRAPH[1499], RIGHT_GRAPH[1435], RIGHT_GRAPH[1371], RIGHT_GRAPH[1307], RIGHT_GRAPH[1243], RIGHT_GRAPH[1179], RIGHT_GRAPH[1115], RIGHT_GRAPH[1051]};
					9'd156	:	PATTERN = {RIGHT_GRAPH[1500], RIGHT_GRAPH[1436], RIGHT_GRAPH[1372], RIGHT_GRAPH[1308], RIGHT_GRAPH[1244], RIGHT_GRAPH[1180], RIGHT_GRAPH[1116], RIGHT_GRAPH[1052]};
					9'd157	:	PATTERN = {RIGHT_GRAPH[1501], RIGHT_GRAPH[1437], RIGHT_GRAPH[1373], RIGHT_GRAPH[1309], RIGHT_GRAPH[1245], RIGHT_GRAPH[1181], RIGHT_GRAPH[1117], RIGHT_GRAPH[1053]};
					9'd158	:	PATTERN = {RIGHT_GRAPH[1502], RIGHT_GRAPH[1438], RIGHT_GRAPH[1374], RIGHT_GRAPH[1310], RIGHT_GRAPH[1246], RIGHT_GRAPH[1182], RIGHT_GRAPH[1118], RIGHT_GRAPH[1054]};
					9'd159	:	PATTERN = {RIGHT_GRAPH[1503], RIGHT_GRAPH[1439], RIGHT_GRAPH[1375], RIGHT_GRAPH[1311], RIGHT_GRAPH[1247], RIGHT_GRAPH[1183], RIGHT_GRAPH[1119], RIGHT_GRAPH[1055]};
					9'd160	:	PATTERN = {RIGHT_GRAPH[1504], RIGHT_GRAPH[1440], RIGHT_GRAPH[1376], RIGHT_GRAPH[1312], RIGHT_GRAPH[1248], RIGHT_GRAPH[1184], RIGHT_GRAPH[1120], RIGHT_GRAPH[1056]};
					9'd161	:	PATTERN = {RIGHT_GRAPH[1505], RIGHT_GRAPH[1441], RIGHT_GRAPH[1377], RIGHT_GRAPH[1313], RIGHT_GRAPH[1249], RIGHT_GRAPH[1185], RIGHT_GRAPH[1121], RIGHT_GRAPH[1057]};
					9'd162	:	PATTERN = {RIGHT_GRAPH[1506], RIGHT_GRAPH[1442], RIGHT_GRAPH[1378], RIGHT_GRAPH[1314], RIGHT_GRAPH[1250], RIGHT_GRAPH[1186], RIGHT_GRAPH[1122], RIGHT_GRAPH[1058]};
					9'd163	:	PATTERN = {RIGHT_GRAPH[1507], RIGHT_GRAPH[1443], RIGHT_GRAPH[1379], RIGHT_GRAPH[1315], RIGHT_GRAPH[1251], RIGHT_GRAPH[1187], RIGHT_GRAPH[1123], RIGHT_GRAPH[1059]};
					9'd164	:	PATTERN = {RIGHT_GRAPH[1508], RIGHT_GRAPH[1444], RIGHT_GRAPH[1380], RIGHT_GRAPH[1316], RIGHT_GRAPH[1252], RIGHT_GRAPH[1188], RIGHT_GRAPH[1124], RIGHT_GRAPH[1060]};
					9'd165	:	PATTERN = {RIGHT_GRAPH[1509], RIGHT_GRAPH[1445], RIGHT_GRAPH[1381], RIGHT_GRAPH[1317], RIGHT_GRAPH[1253], RIGHT_GRAPH[1189], RIGHT_GRAPH[1125], RIGHT_GRAPH[1061]};
					9'd166	:	PATTERN = {RIGHT_GRAPH[1510], RIGHT_GRAPH[1446], RIGHT_GRAPH[1382], RIGHT_GRAPH[1318], RIGHT_GRAPH[1254], RIGHT_GRAPH[1190], RIGHT_GRAPH[1126], RIGHT_GRAPH[1062]};
					9'd167	:	PATTERN = {RIGHT_GRAPH[1511], RIGHT_GRAPH[1447], RIGHT_GRAPH[1383], RIGHT_GRAPH[1319], RIGHT_GRAPH[1255], RIGHT_GRAPH[1191], RIGHT_GRAPH[1127], RIGHT_GRAPH[1063]};
					9'd168	:	PATTERN = {RIGHT_GRAPH[1512], RIGHT_GRAPH[1448], RIGHT_GRAPH[1384], RIGHT_GRAPH[1320], RIGHT_GRAPH[1256], RIGHT_GRAPH[1192], RIGHT_GRAPH[1128], RIGHT_GRAPH[1064]};
					9'd169	:	PATTERN = {RIGHT_GRAPH[1513], RIGHT_GRAPH[1449], RIGHT_GRAPH[1385], RIGHT_GRAPH[1321], RIGHT_GRAPH[1257], RIGHT_GRAPH[1193], RIGHT_GRAPH[1129], RIGHT_GRAPH[1065]};
					9'd170	:	PATTERN = {RIGHT_GRAPH[1514], RIGHT_GRAPH[1450], RIGHT_GRAPH[1386], RIGHT_GRAPH[1322], RIGHT_GRAPH[1258], RIGHT_GRAPH[1194], RIGHT_GRAPH[1130], RIGHT_GRAPH[1066]};
					9'd171	:	PATTERN = {RIGHT_GRAPH[1515], RIGHT_GRAPH[1451], RIGHT_GRAPH[1387], RIGHT_GRAPH[1323], RIGHT_GRAPH[1259], RIGHT_GRAPH[1195], RIGHT_GRAPH[1131], RIGHT_GRAPH[1067]};
					9'd172	:	PATTERN = {RIGHT_GRAPH[1516], RIGHT_GRAPH[1452], RIGHT_GRAPH[1388], RIGHT_GRAPH[1324], RIGHT_GRAPH[1260], RIGHT_GRAPH[1196], RIGHT_GRAPH[1132], RIGHT_GRAPH[1068]};
					9'd173	:	PATTERN = {RIGHT_GRAPH[1517], RIGHT_GRAPH[1453], RIGHT_GRAPH[1389], RIGHT_GRAPH[1325], RIGHT_GRAPH[1261], RIGHT_GRAPH[1197], RIGHT_GRAPH[1133], RIGHT_GRAPH[1069]};
					9'd174	:	PATTERN = {RIGHT_GRAPH[1518], RIGHT_GRAPH[1454], RIGHT_GRAPH[1390], RIGHT_GRAPH[1326], RIGHT_GRAPH[1262], RIGHT_GRAPH[1198], RIGHT_GRAPH[1134], RIGHT_GRAPH[1070]};
					9'd175	:	PATTERN = {RIGHT_GRAPH[1519], RIGHT_GRAPH[1455], RIGHT_GRAPH[1391], RIGHT_GRAPH[1327], RIGHT_GRAPH[1263], RIGHT_GRAPH[1199], RIGHT_GRAPH[1135], RIGHT_GRAPH[1071]};
					9'd176	:	PATTERN = {RIGHT_GRAPH[1520], RIGHT_GRAPH[1456], RIGHT_GRAPH[1392], RIGHT_GRAPH[1328], RIGHT_GRAPH[1264], RIGHT_GRAPH[1200], RIGHT_GRAPH[1136], RIGHT_GRAPH[1072]};
					9'd177	:	PATTERN = {RIGHT_GRAPH[1521], RIGHT_GRAPH[1457], RIGHT_GRAPH[1393], RIGHT_GRAPH[1329], RIGHT_GRAPH[1265], RIGHT_GRAPH[1201], RIGHT_GRAPH[1137], RIGHT_GRAPH[1073]};
					9'd178	:	PATTERN = {RIGHT_GRAPH[1522], RIGHT_GRAPH[1458], RIGHT_GRAPH[1394], RIGHT_GRAPH[1330], RIGHT_GRAPH[1266], RIGHT_GRAPH[1202], RIGHT_GRAPH[1138], RIGHT_GRAPH[1074]};
					9'd179	:	PATTERN = {RIGHT_GRAPH[1523], RIGHT_GRAPH[1459], RIGHT_GRAPH[1395], RIGHT_GRAPH[1331], RIGHT_GRAPH[1267], RIGHT_GRAPH[1203], RIGHT_GRAPH[1139], RIGHT_GRAPH[1075]};
					9'd180	:	PATTERN = {RIGHT_GRAPH[1524], RIGHT_GRAPH[1460], RIGHT_GRAPH[1396], RIGHT_GRAPH[1332], RIGHT_GRAPH[1268], RIGHT_GRAPH[1204], RIGHT_GRAPH[1140], RIGHT_GRAPH[1076]};
					9'd181	:	PATTERN = {RIGHT_GRAPH[1525], RIGHT_GRAPH[1461], RIGHT_GRAPH[1397], RIGHT_GRAPH[1333], RIGHT_GRAPH[1269], RIGHT_GRAPH[1205], RIGHT_GRAPH[1141], RIGHT_GRAPH[1077]};
					9'd182	:	PATTERN = {RIGHT_GRAPH[1526], RIGHT_GRAPH[1462], RIGHT_GRAPH[1398], RIGHT_GRAPH[1334], RIGHT_GRAPH[1270], RIGHT_GRAPH[1206], RIGHT_GRAPH[1142], RIGHT_GRAPH[1078]};
					9'd183	:	PATTERN = {RIGHT_GRAPH[1527], RIGHT_GRAPH[1463], RIGHT_GRAPH[1399], RIGHT_GRAPH[1335], RIGHT_GRAPH[1271], RIGHT_GRAPH[1207], RIGHT_GRAPH[1143], RIGHT_GRAPH[1079]};
					9'd184	:	PATTERN = {RIGHT_GRAPH[1528], RIGHT_GRAPH[1464], RIGHT_GRAPH[1400], RIGHT_GRAPH[1336], RIGHT_GRAPH[1272], RIGHT_GRAPH[1208], RIGHT_GRAPH[1144], RIGHT_GRAPH[1080]};
					9'd185	:	PATTERN = {RIGHT_GRAPH[1529], RIGHT_GRAPH[1465], RIGHT_GRAPH[1401], RIGHT_GRAPH[1337], RIGHT_GRAPH[1273], RIGHT_GRAPH[1209], RIGHT_GRAPH[1145], RIGHT_GRAPH[1081]};
					9'd186	:	PATTERN = {RIGHT_GRAPH[1530], RIGHT_GRAPH[1466], RIGHT_GRAPH[1402], RIGHT_GRAPH[1338], RIGHT_GRAPH[1274], RIGHT_GRAPH[1210], RIGHT_GRAPH[1146], RIGHT_GRAPH[1082]};
					9'd187	:	PATTERN = {RIGHT_GRAPH[1531], RIGHT_GRAPH[1467], RIGHT_GRAPH[1403], RIGHT_GRAPH[1339], RIGHT_GRAPH[1275], RIGHT_GRAPH[1211], RIGHT_GRAPH[1147], RIGHT_GRAPH[1083]};
					9'd188	:	PATTERN = {RIGHT_GRAPH[1532], RIGHT_GRAPH[1468], RIGHT_GRAPH[1404], RIGHT_GRAPH[1340], RIGHT_GRAPH[1276], RIGHT_GRAPH[1212], RIGHT_GRAPH[1148], RIGHT_GRAPH[1084]};
					9'd189	:	PATTERN = {RIGHT_GRAPH[1533], RIGHT_GRAPH[1469], RIGHT_GRAPH[1405], RIGHT_GRAPH[1341], RIGHT_GRAPH[1277], RIGHT_GRAPH[1213], RIGHT_GRAPH[1149], RIGHT_GRAPH[1085]};
					9'd190	:	PATTERN = {RIGHT_GRAPH[1534], RIGHT_GRAPH[1470], RIGHT_GRAPH[1406], RIGHT_GRAPH[1342], RIGHT_GRAPH[1278], RIGHT_GRAPH[1214], RIGHT_GRAPH[1150], RIGHT_GRAPH[1086]};
					9'd191	:	PATTERN = {RIGHT_GRAPH[1535], RIGHT_GRAPH[1471], RIGHT_GRAPH[1407], RIGHT_GRAPH[1343], RIGHT_GRAPH[1279], RIGHT_GRAPH[1215], RIGHT_GRAPH[1151], RIGHT_GRAPH[1087]};
					9'd192	:	PATTERN = {RIGHT_GRAPH[1984], RIGHT_GRAPH[1920], RIGHT_GRAPH[1856], RIGHT_GRAPH[1792], RIGHT_GRAPH[1728], RIGHT_GRAPH[1664], RIGHT_GRAPH[1600], RIGHT_GRAPH[1536]};
					9'd193	:	PATTERN = {RIGHT_GRAPH[1985], RIGHT_GRAPH[1921], RIGHT_GRAPH[1857], RIGHT_GRAPH[1793], RIGHT_GRAPH[1729], RIGHT_GRAPH[1665], RIGHT_GRAPH[1601], RIGHT_GRAPH[1537]};
					9'd194	:	PATTERN = {RIGHT_GRAPH[1986], RIGHT_GRAPH[1922], RIGHT_GRAPH[1858], RIGHT_GRAPH[1794], RIGHT_GRAPH[1730], RIGHT_GRAPH[1666], RIGHT_GRAPH[1602], RIGHT_GRAPH[1538]};
					9'd195	:	PATTERN = {RIGHT_GRAPH[1987], RIGHT_GRAPH[1923], RIGHT_GRAPH[1859], RIGHT_GRAPH[1795], RIGHT_GRAPH[1731], RIGHT_GRAPH[1667], RIGHT_GRAPH[1603], RIGHT_GRAPH[1539]};
					9'd196	:	PATTERN = {RIGHT_GRAPH[1988], RIGHT_GRAPH[1924], RIGHT_GRAPH[1860], RIGHT_GRAPH[1796], RIGHT_GRAPH[1732], RIGHT_GRAPH[1668], RIGHT_GRAPH[1604], RIGHT_GRAPH[1540]};
					9'd197	:	PATTERN = {RIGHT_GRAPH[1989], RIGHT_GRAPH[1925], RIGHT_GRAPH[1861], RIGHT_GRAPH[1797], RIGHT_GRAPH[1733], RIGHT_GRAPH[1669], RIGHT_GRAPH[1605], RIGHT_GRAPH[1541]};
					9'd198	:	PATTERN = {RIGHT_GRAPH[1990], RIGHT_GRAPH[1926], RIGHT_GRAPH[1862], RIGHT_GRAPH[1798], RIGHT_GRAPH[1734], RIGHT_GRAPH[1670], RIGHT_GRAPH[1606], RIGHT_GRAPH[1542]};
					9'd199	:	PATTERN = {RIGHT_GRAPH[1991], RIGHT_GRAPH[1927], RIGHT_GRAPH[1863], RIGHT_GRAPH[1799], RIGHT_GRAPH[1735], RIGHT_GRAPH[1671], RIGHT_GRAPH[1607], RIGHT_GRAPH[1543]};
					9'd200	:	PATTERN = {RIGHT_GRAPH[1992], RIGHT_GRAPH[1928], RIGHT_GRAPH[1864], RIGHT_GRAPH[1800], RIGHT_GRAPH[1736], RIGHT_GRAPH[1672], RIGHT_GRAPH[1608], RIGHT_GRAPH[1544]};
					9'd201	:	PATTERN = {RIGHT_GRAPH[1993], RIGHT_GRAPH[1929], RIGHT_GRAPH[1865], RIGHT_GRAPH[1801], RIGHT_GRAPH[1737], RIGHT_GRAPH[1673], RIGHT_GRAPH[1609], RIGHT_GRAPH[1545]};
					9'd202	:	PATTERN = {RIGHT_GRAPH[1994], RIGHT_GRAPH[1930], RIGHT_GRAPH[1866], RIGHT_GRAPH[1802], RIGHT_GRAPH[1738], RIGHT_GRAPH[1674], RIGHT_GRAPH[1610], RIGHT_GRAPH[1546]};
					9'd203	:	PATTERN = {RIGHT_GRAPH[1995], RIGHT_GRAPH[1931], RIGHT_GRAPH[1867], RIGHT_GRAPH[1803], RIGHT_GRAPH[1739], RIGHT_GRAPH[1675], RIGHT_GRAPH[1611], RIGHT_GRAPH[1547]};
					9'd204	:	PATTERN = {RIGHT_GRAPH[1996], RIGHT_GRAPH[1932], RIGHT_GRAPH[1868], RIGHT_GRAPH[1804], RIGHT_GRAPH[1740], RIGHT_GRAPH[1676], RIGHT_GRAPH[1612], RIGHT_GRAPH[1548]};
					9'd205	:	PATTERN = {RIGHT_GRAPH[1997], RIGHT_GRAPH[1933], RIGHT_GRAPH[1869], RIGHT_GRAPH[1805], RIGHT_GRAPH[1741], RIGHT_GRAPH[1677], RIGHT_GRAPH[1613], RIGHT_GRAPH[1549]};
					9'd206	:	PATTERN = {RIGHT_GRAPH[1998], RIGHT_GRAPH[1934], RIGHT_GRAPH[1870], RIGHT_GRAPH[1806], RIGHT_GRAPH[1742], RIGHT_GRAPH[1678], RIGHT_GRAPH[1614], RIGHT_GRAPH[1550]};
					9'd207	:	PATTERN = {RIGHT_GRAPH[1999], RIGHT_GRAPH[1935], RIGHT_GRAPH[1871], RIGHT_GRAPH[1807], RIGHT_GRAPH[1743], RIGHT_GRAPH[1679], RIGHT_GRAPH[1615], RIGHT_GRAPH[1551]};
					9'd208	:	PATTERN = {RIGHT_GRAPH[2000], RIGHT_GRAPH[1936], RIGHT_GRAPH[1872], RIGHT_GRAPH[1808], RIGHT_GRAPH[1744], RIGHT_GRAPH[1680], RIGHT_GRAPH[1616], RIGHT_GRAPH[1552]};
					9'd209	:	PATTERN = {RIGHT_GRAPH[2001], RIGHT_GRAPH[1937], RIGHT_GRAPH[1873], RIGHT_GRAPH[1809], RIGHT_GRAPH[1745], RIGHT_GRAPH[1681], RIGHT_GRAPH[1617], RIGHT_GRAPH[1553]};
					9'd210	:	PATTERN = {RIGHT_GRAPH[2002], RIGHT_GRAPH[1938], RIGHT_GRAPH[1874], RIGHT_GRAPH[1810], RIGHT_GRAPH[1746], RIGHT_GRAPH[1682], RIGHT_GRAPH[1618], RIGHT_GRAPH[1554]};
					9'd211	:	PATTERN = {RIGHT_GRAPH[2003], RIGHT_GRAPH[1939], RIGHT_GRAPH[1875], RIGHT_GRAPH[1811], RIGHT_GRAPH[1747], RIGHT_GRAPH[1683], RIGHT_GRAPH[1619], RIGHT_GRAPH[1555]};
					9'd212	:	PATTERN = {RIGHT_GRAPH[2004], RIGHT_GRAPH[1940], RIGHT_GRAPH[1876], RIGHT_GRAPH[1812], RIGHT_GRAPH[1748], RIGHT_GRAPH[1684], RIGHT_GRAPH[1620], RIGHT_GRAPH[1556]};
					9'd213	:	PATTERN = {RIGHT_GRAPH[2005], RIGHT_GRAPH[1941], RIGHT_GRAPH[1877], RIGHT_GRAPH[1813], RIGHT_GRAPH[1749], RIGHT_GRAPH[1685], RIGHT_GRAPH[1621], RIGHT_GRAPH[1557]};
					9'd214	:	PATTERN = {RIGHT_GRAPH[2006], RIGHT_GRAPH[1942], RIGHT_GRAPH[1878], RIGHT_GRAPH[1814], RIGHT_GRAPH[1750], RIGHT_GRAPH[1686], RIGHT_GRAPH[1622], RIGHT_GRAPH[1558]};
					9'd215	:	PATTERN = {RIGHT_GRAPH[2007], RIGHT_GRAPH[1943], RIGHT_GRAPH[1879], RIGHT_GRAPH[1815], RIGHT_GRAPH[1751], RIGHT_GRAPH[1687], RIGHT_GRAPH[1623], RIGHT_GRAPH[1559]};
					9'd216	:	PATTERN = {RIGHT_GRAPH[2008], RIGHT_GRAPH[1944], RIGHT_GRAPH[1880], RIGHT_GRAPH[1816], RIGHT_GRAPH[1752], RIGHT_GRAPH[1688], RIGHT_GRAPH[1624], RIGHT_GRAPH[1560]};
					9'd217	:	PATTERN = {RIGHT_GRAPH[2009], RIGHT_GRAPH[1945], RIGHT_GRAPH[1881], RIGHT_GRAPH[1817], RIGHT_GRAPH[1753], RIGHT_GRAPH[1689], RIGHT_GRAPH[1625], RIGHT_GRAPH[1561]};
					9'd218	:	PATTERN = {RIGHT_GRAPH[2010], RIGHT_GRAPH[1946], RIGHT_GRAPH[1882], RIGHT_GRAPH[1818], RIGHT_GRAPH[1754], RIGHT_GRAPH[1690], RIGHT_GRAPH[1626], RIGHT_GRAPH[1562]};
					9'd219	:	PATTERN = {RIGHT_GRAPH[2011], RIGHT_GRAPH[1947], RIGHT_GRAPH[1883], RIGHT_GRAPH[1819], RIGHT_GRAPH[1755], RIGHT_GRAPH[1691], RIGHT_GRAPH[1627], RIGHT_GRAPH[1563]};
					9'd220	:	PATTERN = {RIGHT_GRAPH[2012], RIGHT_GRAPH[1948], RIGHT_GRAPH[1884], RIGHT_GRAPH[1820], RIGHT_GRAPH[1756], RIGHT_GRAPH[1692], RIGHT_GRAPH[1628], RIGHT_GRAPH[1564]};
					9'd221	:	PATTERN = {RIGHT_GRAPH[2013], RIGHT_GRAPH[1949], RIGHT_GRAPH[1885], RIGHT_GRAPH[1821], RIGHT_GRAPH[1757], RIGHT_GRAPH[1693], RIGHT_GRAPH[1629], RIGHT_GRAPH[1565]};
					9'd222	:	PATTERN = {RIGHT_GRAPH[2014], RIGHT_GRAPH[1950], RIGHT_GRAPH[1886], RIGHT_GRAPH[1822], RIGHT_GRAPH[1758], RIGHT_GRAPH[1694], RIGHT_GRAPH[1630], RIGHT_GRAPH[1566]};
					9'd223	:	PATTERN = {RIGHT_GRAPH[2015], RIGHT_GRAPH[1951], RIGHT_GRAPH[1887], RIGHT_GRAPH[1823], RIGHT_GRAPH[1759], RIGHT_GRAPH[1695], RIGHT_GRAPH[1631], RIGHT_GRAPH[1567]};
					9'd224	:	PATTERN = {RIGHT_GRAPH[2016], RIGHT_GRAPH[1952], RIGHT_GRAPH[1888], RIGHT_GRAPH[1824], RIGHT_GRAPH[1760], RIGHT_GRAPH[1696], RIGHT_GRAPH[1632], RIGHT_GRAPH[1568]};
					9'd225	:	PATTERN = {RIGHT_GRAPH[2017], RIGHT_GRAPH[1953], RIGHT_GRAPH[1889], RIGHT_GRAPH[1825], RIGHT_GRAPH[1761], RIGHT_GRAPH[1697], RIGHT_GRAPH[1633], RIGHT_GRAPH[1569]};
					9'd226	:	PATTERN = {RIGHT_GRAPH[2018], RIGHT_GRAPH[1954], RIGHT_GRAPH[1890], RIGHT_GRAPH[1826], RIGHT_GRAPH[1762], RIGHT_GRAPH[1698], RIGHT_GRAPH[1634], RIGHT_GRAPH[1570]};
					9'd227	:	PATTERN = {RIGHT_GRAPH[2019], RIGHT_GRAPH[1955], RIGHT_GRAPH[1891], RIGHT_GRAPH[1827], RIGHT_GRAPH[1763], RIGHT_GRAPH[1699], RIGHT_GRAPH[1635], RIGHT_GRAPH[1571]};
					9'd228	:	PATTERN = {RIGHT_GRAPH[2020], RIGHT_GRAPH[1956], RIGHT_GRAPH[1892], RIGHT_GRAPH[1828], RIGHT_GRAPH[1764], RIGHT_GRAPH[1700], RIGHT_GRAPH[1636], RIGHT_GRAPH[1572]};
					9'd229	:	PATTERN = {RIGHT_GRAPH[2021], RIGHT_GRAPH[1957], RIGHT_GRAPH[1893], RIGHT_GRAPH[1829], RIGHT_GRAPH[1765], RIGHT_GRAPH[1701], RIGHT_GRAPH[1637], RIGHT_GRAPH[1573]};
					9'd230	:	PATTERN = {RIGHT_GRAPH[2022], RIGHT_GRAPH[1958], RIGHT_GRAPH[1894], RIGHT_GRAPH[1830], RIGHT_GRAPH[1766], RIGHT_GRAPH[1702], RIGHT_GRAPH[1638], RIGHT_GRAPH[1574]};
					9'd231	:	PATTERN = {RIGHT_GRAPH[2023], RIGHT_GRAPH[1959], RIGHT_GRAPH[1895], RIGHT_GRAPH[1831], RIGHT_GRAPH[1767], RIGHT_GRAPH[1703], RIGHT_GRAPH[1639], RIGHT_GRAPH[1575]};
					9'd232	:	PATTERN = {RIGHT_GRAPH[2024], RIGHT_GRAPH[1960], RIGHT_GRAPH[1896], RIGHT_GRAPH[1832], RIGHT_GRAPH[1768], RIGHT_GRAPH[1704], RIGHT_GRAPH[1640], RIGHT_GRAPH[1576]};
					9'd233	:	PATTERN = {RIGHT_GRAPH[2025], RIGHT_GRAPH[1961], RIGHT_GRAPH[1897], RIGHT_GRAPH[1833], RIGHT_GRAPH[1769], RIGHT_GRAPH[1705], RIGHT_GRAPH[1641], RIGHT_GRAPH[1577]};
					9'd234	:	PATTERN = {RIGHT_GRAPH[2026], RIGHT_GRAPH[1962], RIGHT_GRAPH[1898], RIGHT_GRAPH[1834], RIGHT_GRAPH[1770], RIGHT_GRAPH[1706], RIGHT_GRAPH[1642], RIGHT_GRAPH[1578]};
					9'd235	:	PATTERN = {RIGHT_GRAPH[2027], RIGHT_GRAPH[1963], RIGHT_GRAPH[1899], RIGHT_GRAPH[1835], RIGHT_GRAPH[1771], RIGHT_GRAPH[1707], RIGHT_GRAPH[1643], RIGHT_GRAPH[1579]};
					9'd236	:	PATTERN = {RIGHT_GRAPH[2028], RIGHT_GRAPH[1964], RIGHT_GRAPH[1900], RIGHT_GRAPH[1836], RIGHT_GRAPH[1772], RIGHT_GRAPH[1708], RIGHT_GRAPH[1644], RIGHT_GRAPH[1580]};
					9'd237	:	PATTERN = {RIGHT_GRAPH[2029], RIGHT_GRAPH[1965], RIGHT_GRAPH[1901], RIGHT_GRAPH[1837], RIGHT_GRAPH[1773], RIGHT_GRAPH[1709], RIGHT_GRAPH[1645], RIGHT_GRAPH[1581]};
					9'd238	:	PATTERN = {RIGHT_GRAPH[2030], RIGHT_GRAPH[1966], RIGHT_GRAPH[1902], RIGHT_GRAPH[1838], RIGHT_GRAPH[1774], RIGHT_GRAPH[1710], RIGHT_GRAPH[1646], RIGHT_GRAPH[1582]};
					9'd239	:	PATTERN = {RIGHT_GRAPH[2031], RIGHT_GRAPH[1967], RIGHT_GRAPH[1903], RIGHT_GRAPH[1839], RIGHT_GRAPH[1775], RIGHT_GRAPH[1711], RIGHT_GRAPH[1647], RIGHT_GRAPH[1583]};
					9'd240	:	PATTERN = {RIGHT_GRAPH[2032], RIGHT_GRAPH[1968], RIGHT_GRAPH[1904], RIGHT_GRAPH[1840], RIGHT_GRAPH[1776], RIGHT_GRAPH[1712], RIGHT_GRAPH[1648], RIGHT_GRAPH[1584]};
					9'd241	:	PATTERN = {RIGHT_GRAPH[2033], RIGHT_GRAPH[1969], RIGHT_GRAPH[1905], RIGHT_GRAPH[1841], RIGHT_GRAPH[1777], RIGHT_GRAPH[1713], RIGHT_GRAPH[1649], RIGHT_GRAPH[1585]};
					9'd242	:	PATTERN = {RIGHT_GRAPH[2034], RIGHT_GRAPH[1970], RIGHT_GRAPH[1906], RIGHT_GRAPH[1842], RIGHT_GRAPH[1778], RIGHT_GRAPH[1714], RIGHT_GRAPH[1650], RIGHT_GRAPH[1586]};
					9'd243	:	PATTERN = {RIGHT_GRAPH[2035], RIGHT_GRAPH[1971], RIGHT_GRAPH[1907], RIGHT_GRAPH[1843], RIGHT_GRAPH[1779], RIGHT_GRAPH[1715], RIGHT_GRAPH[1651], RIGHT_GRAPH[1587]};
					9'd244	:	PATTERN = {RIGHT_GRAPH[2036], RIGHT_GRAPH[1972], RIGHT_GRAPH[1908], RIGHT_GRAPH[1844], RIGHT_GRAPH[1780], RIGHT_GRAPH[1716], RIGHT_GRAPH[1652], RIGHT_GRAPH[1588]};
					9'd245	:	PATTERN = {RIGHT_GRAPH[2037], RIGHT_GRAPH[1973], RIGHT_GRAPH[1909], RIGHT_GRAPH[1845], RIGHT_GRAPH[1781], RIGHT_GRAPH[1717], RIGHT_GRAPH[1653], RIGHT_GRAPH[1589]};
					9'd246	:	PATTERN = {RIGHT_GRAPH[2038], RIGHT_GRAPH[1974], RIGHT_GRAPH[1910], RIGHT_GRAPH[1846], RIGHT_GRAPH[1782], RIGHT_GRAPH[1718], RIGHT_GRAPH[1654], RIGHT_GRAPH[1590]};
					9'd247	:	PATTERN = {RIGHT_GRAPH[2039], RIGHT_GRAPH[1975], RIGHT_GRAPH[1911], RIGHT_GRAPH[1847], RIGHT_GRAPH[1783], RIGHT_GRAPH[1719], RIGHT_GRAPH[1655], RIGHT_GRAPH[1591]};
					9'd248	:	PATTERN = {RIGHT_GRAPH[2040], RIGHT_GRAPH[1976], RIGHT_GRAPH[1912], RIGHT_GRAPH[1848], RIGHT_GRAPH[1784], RIGHT_GRAPH[1720], RIGHT_GRAPH[1656], RIGHT_GRAPH[1592]};
					9'd249	:	PATTERN = {RIGHT_GRAPH[2041], RIGHT_GRAPH[1977], RIGHT_GRAPH[1913], RIGHT_GRAPH[1849], RIGHT_GRAPH[1785], RIGHT_GRAPH[1721], RIGHT_GRAPH[1657], RIGHT_GRAPH[1593]};
					9'd250	:	PATTERN = {RIGHT_GRAPH[2042], RIGHT_GRAPH[1978], RIGHT_GRAPH[1914], RIGHT_GRAPH[1850], RIGHT_GRAPH[1786], RIGHT_GRAPH[1722], RIGHT_GRAPH[1658], RIGHT_GRAPH[1594]};
					9'd251	:	PATTERN = {RIGHT_GRAPH[2043], RIGHT_GRAPH[1979], RIGHT_GRAPH[1915], RIGHT_GRAPH[1851], RIGHT_GRAPH[1787], RIGHT_GRAPH[1723], RIGHT_GRAPH[1659], RIGHT_GRAPH[1595]};
					9'd252	:	PATTERN = {RIGHT_GRAPH[2044], RIGHT_GRAPH[1980], RIGHT_GRAPH[1916], RIGHT_GRAPH[1852], RIGHT_GRAPH[1788], RIGHT_GRAPH[1724], RIGHT_GRAPH[1660], RIGHT_GRAPH[1596]};
					9'd253	:	PATTERN = {RIGHT_GRAPH[2045], RIGHT_GRAPH[1981], RIGHT_GRAPH[1917], RIGHT_GRAPH[1853], RIGHT_GRAPH[1789], RIGHT_GRAPH[1725], RIGHT_GRAPH[1661], RIGHT_GRAPH[1597]};
					9'd254	:	PATTERN = {RIGHT_GRAPH[2046], RIGHT_GRAPH[1982], RIGHT_GRAPH[1918], RIGHT_GRAPH[1854], RIGHT_GRAPH[1790], RIGHT_GRAPH[1726], RIGHT_GRAPH[1662], RIGHT_GRAPH[1598]};
					9'd255	:	PATTERN = {RIGHT_GRAPH[2047], RIGHT_GRAPH[1983], RIGHT_GRAPH[1919], RIGHT_GRAPH[1855], RIGHT_GRAPH[1791], RIGHT_GRAPH[1727], RIGHT_GRAPH[1663], RIGHT_GRAPH[1599]};
					9'd256	:	PATTERN = {RIGHT_GRAPH[2496], RIGHT_GRAPH[2432], RIGHT_GRAPH[2368], RIGHT_GRAPH[2304], RIGHT_GRAPH[2240], RIGHT_GRAPH[2176], RIGHT_GRAPH[2112], RIGHT_GRAPH[2048]};
					9'd257	:	PATTERN = {RIGHT_GRAPH[2497], RIGHT_GRAPH[2433], RIGHT_GRAPH[2369], RIGHT_GRAPH[2305], RIGHT_GRAPH[2241], RIGHT_GRAPH[2177], RIGHT_GRAPH[2113], RIGHT_GRAPH[2049]};
					9'd258	:	PATTERN = {RIGHT_GRAPH[2498], RIGHT_GRAPH[2434], RIGHT_GRAPH[2370], RIGHT_GRAPH[2306], RIGHT_GRAPH[2242], RIGHT_GRAPH[2178], RIGHT_GRAPH[2114], RIGHT_GRAPH[2050]};
					9'd259	:	PATTERN = {RIGHT_GRAPH[2499], RIGHT_GRAPH[2435], RIGHT_GRAPH[2371], RIGHT_GRAPH[2307], RIGHT_GRAPH[2243], RIGHT_GRAPH[2179], RIGHT_GRAPH[2115], RIGHT_GRAPH[2051]};
					9'd260	:	PATTERN = {RIGHT_GRAPH[2500], RIGHT_GRAPH[2436], RIGHT_GRAPH[2372], RIGHT_GRAPH[2308], RIGHT_GRAPH[2244], RIGHT_GRAPH[2180], RIGHT_GRAPH[2116], RIGHT_GRAPH[2052]};
					9'd261	:	PATTERN = {RIGHT_GRAPH[2501], RIGHT_GRAPH[2437], RIGHT_GRAPH[2373], RIGHT_GRAPH[2309], RIGHT_GRAPH[2245], RIGHT_GRAPH[2181], RIGHT_GRAPH[2117], RIGHT_GRAPH[2053]};
					9'd262	:	PATTERN = {RIGHT_GRAPH[2502], RIGHT_GRAPH[2438], RIGHT_GRAPH[2374], RIGHT_GRAPH[2310], RIGHT_GRAPH[2246], RIGHT_GRAPH[2182], RIGHT_GRAPH[2118], RIGHT_GRAPH[2054]};
					9'd263	:	PATTERN = {RIGHT_GRAPH[2503], RIGHT_GRAPH[2439], RIGHT_GRAPH[2375], RIGHT_GRAPH[2311], RIGHT_GRAPH[2247], RIGHT_GRAPH[2183], RIGHT_GRAPH[2119], RIGHT_GRAPH[2055]};
					9'd264	:	PATTERN = {RIGHT_GRAPH[2504], RIGHT_GRAPH[2440], RIGHT_GRAPH[2376], RIGHT_GRAPH[2312], RIGHT_GRAPH[2248], RIGHT_GRAPH[2184], RIGHT_GRAPH[2120], RIGHT_GRAPH[2056]};
					9'd265	:	PATTERN = {RIGHT_GRAPH[2505], RIGHT_GRAPH[2441], RIGHT_GRAPH[2377], RIGHT_GRAPH[2313], RIGHT_GRAPH[2249], RIGHT_GRAPH[2185], RIGHT_GRAPH[2121], RIGHT_GRAPH[2057]};
					9'd266	:	PATTERN = {RIGHT_GRAPH[2506], RIGHT_GRAPH[2442], RIGHT_GRAPH[2378], RIGHT_GRAPH[2314], RIGHT_GRAPH[2250], RIGHT_GRAPH[2186], RIGHT_GRAPH[2122], RIGHT_GRAPH[2058]};
					9'd267	:	PATTERN = {RIGHT_GRAPH[2507], RIGHT_GRAPH[2443], RIGHT_GRAPH[2379], RIGHT_GRAPH[2315], RIGHT_GRAPH[2251], RIGHT_GRAPH[2187], RIGHT_GRAPH[2123], RIGHT_GRAPH[2059]};
					9'd268	:	PATTERN = {RIGHT_GRAPH[2508], RIGHT_GRAPH[2444], RIGHT_GRAPH[2380], RIGHT_GRAPH[2316], RIGHT_GRAPH[2252], RIGHT_GRAPH[2188], RIGHT_GRAPH[2124], RIGHT_GRAPH[2060]};
					9'd269	:	PATTERN = {RIGHT_GRAPH[2509], RIGHT_GRAPH[2445], RIGHT_GRAPH[2381], RIGHT_GRAPH[2317], RIGHT_GRAPH[2253], RIGHT_GRAPH[2189], RIGHT_GRAPH[2125], RIGHT_GRAPH[2061]};
					9'd270	:	PATTERN = {RIGHT_GRAPH[2510], RIGHT_GRAPH[2446], RIGHT_GRAPH[2382], RIGHT_GRAPH[2318], RIGHT_GRAPH[2254], RIGHT_GRAPH[2190], RIGHT_GRAPH[2126], RIGHT_GRAPH[2062]};
					9'd271	:	PATTERN = {RIGHT_GRAPH[2511], RIGHT_GRAPH[2447], RIGHT_GRAPH[2383], RIGHT_GRAPH[2319], RIGHT_GRAPH[2255], RIGHT_GRAPH[2191], RIGHT_GRAPH[2127], RIGHT_GRAPH[2063]};
					9'd272	:	PATTERN = {RIGHT_GRAPH[2512], RIGHT_GRAPH[2448], RIGHT_GRAPH[2384], RIGHT_GRAPH[2320], RIGHT_GRAPH[2256], RIGHT_GRAPH[2192], RIGHT_GRAPH[2128], RIGHT_GRAPH[2064]};
					9'd273	:	PATTERN = {RIGHT_GRAPH[2513], RIGHT_GRAPH[2449], RIGHT_GRAPH[2385], RIGHT_GRAPH[2321], RIGHT_GRAPH[2257], RIGHT_GRAPH[2193], RIGHT_GRAPH[2129], RIGHT_GRAPH[2065]};
					9'd274	:	PATTERN = {RIGHT_GRAPH[2514], RIGHT_GRAPH[2450], RIGHT_GRAPH[2386], RIGHT_GRAPH[2322], RIGHT_GRAPH[2258], RIGHT_GRAPH[2194], RIGHT_GRAPH[2130], RIGHT_GRAPH[2066]};
					9'd275	:	PATTERN = {RIGHT_GRAPH[2515], RIGHT_GRAPH[2451], RIGHT_GRAPH[2387], RIGHT_GRAPH[2323], RIGHT_GRAPH[2259], RIGHT_GRAPH[2195], RIGHT_GRAPH[2131], RIGHT_GRAPH[2067]};
					9'd276	:	PATTERN = {RIGHT_GRAPH[2516], RIGHT_GRAPH[2452], RIGHT_GRAPH[2388], RIGHT_GRAPH[2324], RIGHT_GRAPH[2260], RIGHT_GRAPH[2196], RIGHT_GRAPH[2132], RIGHT_GRAPH[2068]};
					9'd277	:	PATTERN = {RIGHT_GRAPH[2517], RIGHT_GRAPH[2453], RIGHT_GRAPH[2389], RIGHT_GRAPH[2325], RIGHT_GRAPH[2261], RIGHT_GRAPH[2197], RIGHT_GRAPH[2133], RIGHT_GRAPH[2069]};
					9'd278	:	PATTERN = {RIGHT_GRAPH[2518], RIGHT_GRAPH[2454], RIGHT_GRAPH[2390], RIGHT_GRAPH[2326], RIGHT_GRAPH[2262], RIGHT_GRAPH[2198], RIGHT_GRAPH[2134], RIGHT_GRAPH[2070]};
					9'd279	:	PATTERN = {RIGHT_GRAPH[2519], RIGHT_GRAPH[2455], RIGHT_GRAPH[2391], RIGHT_GRAPH[2327], RIGHT_GRAPH[2263], RIGHT_GRAPH[2199], RIGHT_GRAPH[2135], RIGHT_GRAPH[2071]};
					9'd280	:	PATTERN = {RIGHT_GRAPH[2520], RIGHT_GRAPH[2456], RIGHT_GRAPH[2392], RIGHT_GRAPH[2328], RIGHT_GRAPH[2264], RIGHT_GRAPH[2200], RIGHT_GRAPH[2136], RIGHT_GRAPH[2072]};
					9'd281	:	PATTERN = {RIGHT_GRAPH[2521], RIGHT_GRAPH[2457], RIGHT_GRAPH[2393], RIGHT_GRAPH[2329], RIGHT_GRAPH[2265], RIGHT_GRAPH[2201], RIGHT_GRAPH[2137], RIGHT_GRAPH[2073]};
					9'd282	:	PATTERN = {RIGHT_GRAPH[2522], RIGHT_GRAPH[2458], RIGHT_GRAPH[2394], RIGHT_GRAPH[2330], RIGHT_GRAPH[2266], RIGHT_GRAPH[2202], RIGHT_GRAPH[2138], RIGHT_GRAPH[2074]};
					9'd283	:	PATTERN = {RIGHT_GRAPH[2523], RIGHT_GRAPH[2459], RIGHT_GRAPH[2395], RIGHT_GRAPH[2331], RIGHT_GRAPH[2267], RIGHT_GRAPH[2203], RIGHT_GRAPH[2139], RIGHT_GRAPH[2075]};
					9'd284	:	PATTERN = {RIGHT_GRAPH[2524], RIGHT_GRAPH[2460], RIGHT_GRAPH[2396], RIGHT_GRAPH[2332], RIGHT_GRAPH[2268], RIGHT_GRAPH[2204], RIGHT_GRAPH[2140], RIGHT_GRAPH[2076]};
					9'd285	:	PATTERN = {RIGHT_GRAPH[2525], RIGHT_GRAPH[2461], RIGHT_GRAPH[2397], RIGHT_GRAPH[2333], RIGHT_GRAPH[2269], RIGHT_GRAPH[2205], RIGHT_GRAPH[2141], RIGHT_GRAPH[2077]};
					9'd286	:	PATTERN = {RIGHT_GRAPH[2526], RIGHT_GRAPH[2462], RIGHT_GRAPH[2398], RIGHT_GRAPH[2334], RIGHT_GRAPH[2270], RIGHT_GRAPH[2206], RIGHT_GRAPH[2142], RIGHT_GRAPH[2078]};
					9'd287	:	PATTERN = {RIGHT_GRAPH[2527], RIGHT_GRAPH[2463], RIGHT_GRAPH[2399], RIGHT_GRAPH[2335], RIGHT_GRAPH[2271], RIGHT_GRAPH[2207], RIGHT_GRAPH[2143], RIGHT_GRAPH[2079]};
					9'd288	:	PATTERN = {RIGHT_GRAPH[2528], RIGHT_GRAPH[2464], RIGHT_GRAPH[2400], RIGHT_GRAPH[2336], RIGHT_GRAPH[2272], RIGHT_GRAPH[2208], RIGHT_GRAPH[2144], RIGHT_GRAPH[2080]};
					9'd289	:	PATTERN = {RIGHT_GRAPH[2529], RIGHT_GRAPH[2465], RIGHT_GRAPH[2401], RIGHT_GRAPH[2337], RIGHT_GRAPH[2273], RIGHT_GRAPH[2209], RIGHT_GRAPH[2145], RIGHT_GRAPH[2081]};
					9'd290	:	PATTERN = {RIGHT_GRAPH[2530], RIGHT_GRAPH[2466], RIGHT_GRAPH[2402], RIGHT_GRAPH[2338], RIGHT_GRAPH[2274], RIGHT_GRAPH[2210], RIGHT_GRAPH[2146], RIGHT_GRAPH[2082]};
					9'd291	:	PATTERN = {RIGHT_GRAPH[2531], RIGHT_GRAPH[2467], RIGHT_GRAPH[2403], RIGHT_GRAPH[2339], RIGHT_GRAPH[2275], RIGHT_GRAPH[2211], RIGHT_GRAPH[2147], RIGHT_GRAPH[2083]};
					9'd292	:	PATTERN = {RIGHT_GRAPH[2532], RIGHT_GRAPH[2468], RIGHT_GRAPH[2404], RIGHT_GRAPH[2340], RIGHT_GRAPH[2276], RIGHT_GRAPH[2212], RIGHT_GRAPH[2148], RIGHT_GRAPH[2084]};
					9'd293	:	PATTERN = {RIGHT_GRAPH[2533], RIGHT_GRAPH[2469], RIGHT_GRAPH[2405], RIGHT_GRAPH[2341], RIGHT_GRAPH[2277], RIGHT_GRAPH[2213], RIGHT_GRAPH[2149], RIGHT_GRAPH[2085]};
					9'd294	:	PATTERN = {RIGHT_GRAPH[2534], RIGHT_GRAPH[2470], RIGHT_GRAPH[2406], RIGHT_GRAPH[2342], RIGHT_GRAPH[2278], RIGHT_GRAPH[2214], RIGHT_GRAPH[2150], RIGHT_GRAPH[2086]};
					9'd295	:	PATTERN = {RIGHT_GRAPH[2535], RIGHT_GRAPH[2471], RIGHT_GRAPH[2407], RIGHT_GRAPH[2343], RIGHT_GRAPH[2279], RIGHT_GRAPH[2215], RIGHT_GRAPH[2151], RIGHT_GRAPH[2087]};
					9'd296	:	PATTERN = {RIGHT_GRAPH[2536], RIGHT_GRAPH[2472], RIGHT_GRAPH[2408], RIGHT_GRAPH[2344], RIGHT_GRAPH[2280], RIGHT_GRAPH[2216], RIGHT_GRAPH[2152], RIGHT_GRAPH[2088]};
					9'd297	:	PATTERN = {RIGHT_GRAPH[2537], RIGHT_GRAPH[2473], RIGHT_GRAPH[2409], RIGHT_GRAPH[2345], RIGHT_GRAPH[2281], RIGHT_GRAPH[2217], RIGHT_GRAPH[2153], RIGHT_GRAPH[2089]};
					9'd298	:	PATTERN = {RIGHT_GRAPH[2538], RIGHT_GRAPH[2474], RIGHT_GRAPH[2410], RIGHT_GRAPH[2346], RIGHT_GRAPH[2282], RIGHT_GRAPH[2218], RIGHT_GRAPH[2154], RIGHT_GRAPH[2090]};
					9'd299	:	PATTERN = {RIGHT_GRAPH[2539], RIGHT_GRAPH[2475], RIGHT_GRAPH[2411], RIGHT_GRAPH[2347], RIGHT_GRAPH[2283], RIGHT_GRAPH[2219], RIGHT_GRAPH[2155], RIGHT_GRAPH[2091]};
					9'd300	:	PATTERN = {RIGHT_GRAPH[2540], RIGHT_GRAPH[2476], RIGHT_GRAPH[2412], RIGHT_GRAPH[2348], RIGHT_GRAPH[2284], RIGHT_GRAPH[2220], RIGHT_GRAPH[2156], RIGHT_GRAPH[2092]};
					9'd301	:	PATTERN = {RIGHT_GRAPH[2541], RIGHT_GRAPH[2477], RIGHT_GRAPH[2413], RIGHT_GRAPH[2349], RIGHT_GRAPH[2285], RIGHT_GRAPH[2221], RIGHT_GRAPH[2157], RIGHT_GRAPH[2093]};
					9'd302	:	PATTERN = {RIGHT_GRAPH[2542], RIGHT_GRAPH[2478], RIGHT_GRAPH[2414], RIGHT_GRAPH[2350], RIGHT_GRAPH[2286], RIGHT_GRAPH[2222], RIGHT_GRAPH[2158], RIGHT_GRAPH[2094]};
					9'd303	:	PATTERN = {RIGHT_GRAPH[2543], RIGHT_GRAPH[2479], RIGHT_GRAPH[2415], RIGHT_GRAPH[2351], RIGHT_GRAPH[2287], RIGHT_GRAPH[2223], RIGHT_GRAPH[2159], RIGHT_GRAPH[2095]};
					9'd304	:	PATTERN = {RIGHT_GRAPH[2544], RIGHT_GRAPH[2480], RIGHT_GRAPH[2416], RIGHT_GRAPH[2352], RIGHT_GRAPH[2288], RIGHT_GRAPH[2224], RIGHT_GRAPH[2160], RIGHT_GRAPH[2096]};
					9'd305	:	PATTERN = {RIGHT_GRAPH[2545], RIGHT_GRAPH[2481], RIGHT_GRAPH[2417], RIGHT_GRAPH[2353], RIGHT_GRAPH[2289], RIGHT_GRAPH[2225], RIGHT_GRAPH[2161], RIGHT_GRAPH[2097]};
					9'd306	:	PATTERN = {RIGHT_GRAPH[2546], RIGHT_GRAPH[2482], RIGHT_GRAPH[2418], RIGHT_GRAPH[2354], RIGHT_GRAPH[2290], RIGHT_GRAPH[2226], RIGHT_GRAPH[2162], RIGHT_GRAPH[2098]};
					9'd307	:	PATTERN = {RIGHT_GRAPH[2547], RIGHT_GRAPH[2483], RIGHT_GRAPH[2419], RIGHT_GRAPH[2355], RIGHT_GRAPH[2291], RIGHT_GRAPH[2227], RIGHT_GRAPH[2163], RIGHT_GRAPH[2099]};
					9'd308	:	PATTERN = {RIGHT_GRAPH[2548], RIGHT_GRAPH[2484], RIGHT_GRAPH[2420], RIGHT_GRAPH[2356], RIGHT_GRAPH[2292], RIGHT_GRAPH[2228], RIGHT_GRAPH[2164], RIGHT_GRAPH[2100]};
					9'd309	:	PATTERN = {RIGHT_GRAPH[2549], RIGHT_GRAPH[2485], RIGHT_GRAPH[2421], RIGHT_GRAPH[2357], RIGHT_GRAPH[2293], RIGHT_GRAPH[2229], RIGHT_GRAPH[2165], RIGHT_GRAPH[2101]};
					9'd310	:	PATTERN = {RIGHT_GRAPH[2550], RIGHT_GRAPH[2486], RIGHT_GRAPH[2422], RIGHT_GRAPH[2358], RIGHT_GRAPH[2294], RIGHT_GRAPH[2230], RIGHT_GRAPH[2166], RIGHT_GRAPH[2102]};
					9'd311	:	PATTERN = {RIGHT_GRAPH[2551], RIGHT_GRAPH[2487], RIGHT_GRAPH[2423], RIGHT_GRAPH[2359], RIGHT_GRAPH[2295], RIGHT_GRAPH[2231], RIGHT_GRAPH[2167], RIGHT_GRAPH[2103]};
					9'd312	:	PATTERN = {RIGHT_GRAPH[2552], RIGHT_GRAPH[2488], RIGHT_GRAPH[2424], RIGHT_GRAPH[2360], RIGHT_GRAPH[2296], RIGHT_GRAPH[2232], RIGHT_GRAPH[2168], RIGHT_GRAPH[2104]};
					9'd313	:	PATTERN = {RIGHT_GRAPH[2553], RIGHT_GRAPH[2489], RIGHT_GRAPH[2425], RIGHT_GRAPH[2361], RIGHT_GRAPH[2297], RIGHT_GRAPH[2233], RIGHT_GRAPH[2169], RIGHT_GRAPH[2105]};
					9'd314	:	PATTERN = {RIGHT_GRAPH[2554], RIGHT_GRAPH[2490], RIGHT_GRAPH[2426], RIGHT_GRAPH[2362], RIGHT_GRAPH[2298], RIGHT_GRAPH[2234], RIGHT_GRAPH[2170], RIGHT_GRAPH[2106]};
					9'd315	:	PATTERN = {RIGHT_GRAPH[2555], RIGHT_GRAPH[2491], RIGHT_GRAPH[2427], RIGHT_GRAPH[2363], RIGHT_GRAPH[2299], RIGHT_GRAPH[2235], RIGHT_GRAPH[2171], RIGHT_GRAPH[2107]};
					9'd316	:	PATTERN = {RIGHT_GRAPH[2556], RIGHT_GRAPH[2492], RIGHT_GRAPH[2428], RIGHT_GRAPH[2364], RIGHT_GRAPH[2300], RIGHT_GRAPH[2236], RIGHT_GRAPH[2172], RIGHT_GRAPH[2108]};
					9'd317	:	PATTERN = {RIGHT_GRAPH[2557], RIGHT_GRAPH[2493], RIGHT_GRAPH[2429], RIGHT_GRAPH[2365], RIGHT_GRAPH[2301], RIGHT_GRAPH[2237], RIGHT_GRAPH[2173], RIGHT_GRAPH[2109]};
					9'd318	:	PATTERN = {RIGHT_GRAPH[2558], RIGHT_GRAPH[2494], RIGHT_GRAPH[2430], RIGHT_GRAPH[2366], RIGHT_GRAPH[2302], RIGHT_GRAPH[2238], RIGHT_GRAPH[2174], RIGHT_GRAPH[2110]};
					9'd319	:	PATTERN = {RIGHT_GRAPH[2559], RIGHT_GRAPH[2495], RIGHT_GRAPH[2431], RIGHT_GRAPH[2367], RIGHT_GRAPH[2303], RIGHT_GRAPH[2239], RIGHT_GRAPH[2175], RIGHT_GRAPH[2111]};
					9'd320	:	PATTERN = {RIGHT_GRAPH[3008], RIGHT_GRAPH[2944], RIGHT_GRAPH[2880], RIGHT_GRAPH[2816], RIGHT_GRAPH[2752], RIGHT_GRAPH[2688], RIGHT_GRAPH[2624], RIGHT_GRAPH[2560]};
					9'd321	:	PATTERN = {RIGHT_GRAPH[3009], RIGHT_GRAPH[2945], RIGHT_GRAPH[2881], RIGHT_GRAPH[2817], RIGHT_GRAPH[2753], RIGHT_GRAPH[2689], RIGHT_GRAPH[2625], RIGHT_GRAPH[2561]};
					9'd322	:	PATTERN = {RIGHT_GRAPH[3010], RIGHT_GRAPH[2946], RIGHT_GRAPH[2882], RIGHT_GRAPH[2818], RIGHT_GRAPH[2754], RIGHT_GRAPH[2690], RIGHT_GRAPH[2626], RIGHT_GRAPH[2562]};
					9'd323	:	PATTERN = {RIGHT_GRAPH[3011], RIGHT_GRAPH[2947], RIGHT_GRAPH[2883], RIGHT_GRAPH[2819], RIGHT_GRAPH[2755], RIGHT_GRAPH[2691], RIGHT_GRAPH[2627], RIGHT_GRAPH[2563]};
					9'd324	:	PATTERN = {RIGHT_GRAPH[3012], RIGHT_GRAPH[2948], RIGHT_GRAPH[2884], RIGHT_GRAPH[2820], RIGHT_GRAPH[2756], RIGHT_GRAPH[2692], RIGHT_GRAPH[2628], RIGHT_GRAPH[2564]};
					9'd325	:	PATTERN = {RIGHT_GRAPH[3013], RIGHT_GRAPH[2949], RIGHT_GRAPH[2885], RIGHT_GRAPH[2821], RIGHT_GRAPH[2757], RIGHT_GRAPH[2693], RIGHT_GRAPH[2629], RIGHT_GRAPH[2565]};
					9'd326	:	PATTERN = {RIGHT_GRAPH[3014], RIGHT_GRAPH[2950], RIGHT_GRAPH[2886], RIGHT_GRAPH[2822], RIGHT_GRAPH[2758], RIGHT_GRAPH[2694], RIGHT_GRAPH[2630], RIGHT_GRAPH[2566]};
					9'd327	:	PATTERN = {RIGHT_GRAPH[3015], RIGHT_GRAPH[2951], RIGHT_GRAPH[2887], RIGHT_GRAPH[2823], RIGHT_GRAPH[2759], RIGHT_GRAPH[2695], RIGHT_GRAPH[2631], RIGHT_GRAPH[2567]};
					9'd328	:	PATTERN = {RIGHT_GRAPH[3016], RIGHT_GRAPH[2952], RIGHT_GRAPH[2888], RIGHT_GRAPH[2824], RIGHT_GRAPH[2760], RIGHT_GRAPH[2696], RIGHT_GRAPH[2632], RIGHT_GRAPH[2568]};
					9'd329	:	PATTERN = {RIGHT_GRAPH[3017], RIGHT_GRAPH[2953], RIGHT_GRAPH[2889], RIGHT_GRAPH[2825], RIGHT_GRAPH[2761], RIGHT_GRAPH[2697], RIGHT_GRAPH[2633], RIGHT_GRAPH[2569]};
					9'd330	:	PATTERN = {RIGHT_GRAPH[3018], RIGHT_GRAPH[2954], RIGHT_GRAPH[2890], RIGHT_GRAPH[2826], RIGHT_GRAPH[2762], RIGHT_GRAPH[2698], RIGHT_GRAPH[2634], RIGHT_GRAPH[2570]};
					9'd331	:	PATTERN = {RIGHT_GRAPH[3019], RIGHT_GRAPH[2955], RIGHT_GRAPH[2891], RIGHT_GRAPH[2827], RIGHT_GRAPH[2763], RIGHT_GRAPH[2699], RIGHT_GRAPH[2635], RIGHT_GRAPH[2571]};
					9'd332	:	PATTERN = {RIGHT_GRAPH[3020], RIGHT_GRAPH[2956], RIGHT_GRAPH[2892], RIGHT_GRAPH[2828], RIGHT_GRAPH[2764], RIGHT_GRAPH[2700], RIGHT_GRAPH[2636], RIGHT_GRAPH[2572]};
					9'd333	:	PATTERN = {RIGHT_GRAPH[3021], RIGHT_GRAPH[2957], RIGHT_GRAPH[2893], RIGHT_GRAPH[2829], RIGHT_GRAPH[2765], RIGHT_GRAPH[2701], RIGHT_GRAPH[2637], RIGHT_GRAPH[2573]};
					9'd334	:	PATTERN = {RIGHT_GRAPH[3022], RIGHT_GRAPH[2958], RIGHT_GRAPH[2894], RIGHT_GRAPH[2830], RIGHT_GRAPH[2766], RIGHT_GRAPH[2702], RIGHT_GRAPH[2638], RIGHT_GRAPH[2574]};
					9'd335	:	PATTERN = {RIGHT_GRAPH[3023], RIGHT_GRAPH[2959], RIGHT_GRAPH[2895], RIGHT_GRAPH[2831], RIGHT_GRAPH[2767], RIGHT_GRAPH[2703], RIGHT_GRAPH[2639], RIGHT_GRAPH[2575]};
					9'd336	:	PATTERN = {RIGHT_GRAPH[3024], RIGHT_GRAPH[2960], RIGHT_GRAPH[2896], RIGHT_GRAPH[2832], RIGHT_GRAPH[2768], RIGHT_GRAPH[2704], RIGHT_GRAPH[2640], RIGHT_GRAPH[2576]};
					9'd337	:	PATTERN = {RIGHT_GRAPH[3025], RIGHT_GRAPH[2961], RIGHT_GRAPH[2897], RIGHT_GRAPH[2833], RIGHT_GRAPH[2769], RIGHT_GRAPH[2705], RIGHT_GRAPH[2641], RIGHT_GRAPH[2577]};
					9'd338	:	PATTERN = {RIGHT_GRAPH[3026], RIGHT_GRAPH[2962], RIGHT_GRAPH[2898], RIGHT_GRAPH[2834], RIGHT_GRAPH[2770], RIGHT_GRAPH[2706], RIGHT_GRAPH[2642], RIGHT_GRAPH[2578]};
					9'd339	:	PATTERN = {RIGHT_GRAPH[3027], RIGHT_GRAPH[2963], RIGHT_GRAPH[2899], RIGHT_GRAPH[2835], RIGHT_GRAPH[2771], RIGHT_GRAPH[2707], RIGHT_GRAPH[2643], RIGHT_GRAPH[2579]};
					9'd340	:	PATTERN = {RIGHT_GRAPH[3028], RIGHT_GRAPH[2964], RIGHT_GRAPH[2900], RIGHT_GRAPH[2836], RIGHT_GRAPH[2772], RIGHT_GRAPH[2708], RIGHT_GRAPH[2644], RIGHT_GRAPH[2580]};
					9'd341	:	PATTERN = {RIGHT_GRAPH[3029], RIGHT_GRAPH[2965], RIGHT_GRAPH[2901], RIGHT_GRAPH[2837], RIGHT_GRAPH[2773], RIGHT_GRAPH[2709], RIGHT_GRAPH[2645], RIGHT_GRAPH[2581]};
					9'd342	:	PATTERN = {RIGHT_GRAPH[3030], RIGHT_GRAPH[2966], RIGHT_GRAPH[2902], RIGHT_GRAPH[2838], RIGHT_GRAPH[2774], RIGHT_GRAPH[2710], RIGHT_GRAPH[2646], RIGHT_GRAPH[2582]};
					9'd343	:	PATTERN = {RIGHT_GRAPH[3031], RIGHT_GRAPH[2967], RIGHT_GRAPH[2903], RIGHT_GRAPH[2839], RIGHT_GRAPH[2775], RIGHT_GRAPH[2711], RIGHT_GRAPH[2647], RIGHT_GRAPH[2583]};
					9'd344	:	PATTERN = {RIGHT_GRAPH[3032], RIGHT_GRAPH[2968], RIGHT_GRAPH[2904], RIGHT_GRAPH[2840], RIGHT_GRAPH[2776], RIGHT_GRAPH[2712], RIGHT_GRAPH[2648], RIGHT_GRAPH[2584]};
					9'd345	:	PATTERN = {RIGHT_GRAPH[3033], RIGHT_GRAPH[2969], RIGHT_GRAPH[2905], RIGHT_GRAPH[2841], RIGHT_GRAPH[2777], RIGHT_GRAPH[2713], RIGHT_GRAPH[2649], RIGHT_GRAPH[2585]};
					9'd346	:	PATTERN = {RIGHT_GRAPH[3034], RIGHT_GRAPH[2970], RIGHT_GRAPH[2906], RIGHT_GRAPH[2842], RIGHT_GRAPH[2778], RIGHT_GRAPH[2714], RIGHT_GRAPH[2650], RIGHT_GRAPH[2586]};
					9'd347	:	PATTERN = {RIGHT_GRAPH[3035], RIGHT_GRAPH[2971], RIGHT_GRAPH[2907], RIGHT_GRAPH[2843], RIGHT_GRAPH[2779], RIGHT_GRAPH[2715], RIGHT_GRAPH[2651], RIGHT_GRAPH[2587]};
					9'd348	:	PATTERN = {RIGHT_GRAPH[3036], RIGHT_GRAPH[2972], RIGHT_GRAPH[2908], RIGHT_GRAPH[2844], RIGHT_GRAPH[2780], RIGHT_GRAPH[2716], RIGHT_GRAPH[2652], RIGHT_GRAPH[2588]};
					9'd349	:	PATTERN = {RIGHT_GRAPH[3037], RIGHT_GRAPH[2973], RIGHT_GRAPH[2909], RIGHT_GRAPH[2845], RIGHT_GRAPH[2781], RIGHT_GRAPH[2717], RIGHT_GRAPH[2653], RIGHT_GRAPH[2589]};
					9'd350	:	PATTERN = {RIGHT_GRAPH[3038], RIGHT_GRAPH[2974], RIGHT_GRAPH[2910], RIGHT_GRAPH[2846], RIGHT_GRAPH[2782], RIGHT_GRAPH[2718], RIGHT_GRAPH[2654], RIGHT_GRAPH[2590]};
					9'd351	:	PATTERN = {RIGHT_GRAPH[3039], RIGHT_GRAPH[2975], RIGHT_GRAPH[2911], RIGHT_GRAPH[2847], RIGHT_GRAPH[2783], RIGHT_GRAPH[2719], RIGHT_GRAPH[2655], RIGHT_GRAPH[2591]};
					9'd352	:	PATTERN = {RIGHT_GRAPH[3040], RIGHT_GRAPH[2976], RIGHT_GRAPH[2912], RIGHT_GRAPH[2848], RIGHT_GRAPH[2784], RIGHT_GRAPH[2720], RIGHT_GRAPH[2656], RIGHT_GRAPH[2592]};
					9'd353	:	PATTERN = {RIGHT_GRAPH[3041], RIGHT_GRAPH[2977], RIGHT_GRAPH[2913], RIGHT_GRAPH[2849], RIGHT_GRAPH[2785], RIGHT_GRAPH[2721], RIGHT_GRAPH[2657], RIGHT_GRAPH[2593]};
					9'd354	:	PATTERN = {RIGHT_GRAPH[3042], RIGHT_GRAPH[2978], RIGHT_GRAPH[2914], RIGHT_GRAPH[2850], RIGHT_GRAPH[2786], RIGHT_GRAPH[2722], RIGHT_GRAPH[2658], RIGHT_GRAPH[2594]};
					9'd355	:	PATTERN = {RIGHT_GRAPH[3043], RIGHT_GRAPH[2979], RIGHT_GRAPH[2915], RIGHT_GRAPH[2851], RIGHT_GRAPH[2787], RIGHT_GRAPH[2723], RIGHT_GRAPH[2659], RIGHT_GRAPH[2595]};
					9'd356	:	PATTERN = {RIGHT_GRAPH[3044], RIGHT_GRAPH[2980], RIGHT_GRAPH[2916], RIGHT_GRAPH[2852], RIGHT_GRAPH[2788], RIGHT_GRAPH[2724], RIGHT_GRAPH[2660], RIGHT_GRAPH[2596]};
					9'd357	:	PATTERN = {RIGHT_GRAPH[3045], RIGHT_GRAPH[2981], RIGHT_GRAPH[2917], RIGHT_GRAPH[2853], RIGHT_GRAPH[2789], RIGHT_GRAPH[2725], RIGHT_GRAPH[2661], RIGHT_GRAPH[2597]};
					9'd358	:	PATTERN = {RIGHT_GRAPH[3046], RIGHT_GRAPH[2982], RIGHT_GRAPH[2918], RIGHT_GRAPH[2854], RIGHT_GRAPH[2790], RIGHT_GRAPH[2726], RIGHT_GRAPH[2662], RIGHT_GRAPH[2598]};
					9'd359	:	PATTERN = {RIGHT_GRAPH[3047], RIGHT_GRAPH[2983], RIGHT_GRAPH[2919], RIGHT_GRAPH[2855], RIGHT_GRAPH[2791], RIGHT_GRAPH[2727], RIGHT_GRAPH[2663], RIGHT_GRAPH[2599]};
					9'd360	:	PATTERN = {RIGHT_GRAPH[3048], RIGHT_GRAPH[2984], RIGHT_GRAPH[2920], RIGHT_GRAPH[2856], RIGHT_GRAPH[2792], RIGHT_GRAPH[2728], RIGHT_GRAPH[2664], RIGHT_GRAPH[2600]};
					9'd361	:	PATTERN = {RIGHT_GRAPH[3049], RIGHT_GRAPH[2985], RIGHT_GRAPH[2921], RIGHT_GRAPH[2857], RIGHT_GRAPH[2793], RIGHT_GRAPH[2729], RIGHT_GRAPH[2665], RIGHT_GRAPH[2601]};
					9'd362	:	PATTERN = {RIGHT_GRAPH[3050], RIGHT_GRAPH[2986], RIGHT_GRAPH[2922], RIGHT_GRAPH[2858], RIGHT_GRAPH[2794], RIGHT_GRAPH[2730], RIGHT_GRAPH[2666], RIGHT_GRAPH[2602]};
					9'd363	:	PATTERN = {RIGHT_GRAPH[3051], RIGHT_GRAPH[2987], RIGHT_GRAPH[2923], RIGHT_GRAPH[2859], RIGHT_GRAPH[2795], RIGHT_GRAPH[2731], RIGHT_GRAPH[2667], RIGHT_GRAPH[2603]};
					9'd364	:	PATTERN = {RIGHT_GRAPH[3052], RIGHT_GRAPH[2988], RIGHT_GRAPH[2924], RIGHT_GRAPH[2860], RIGHT_GRAPH[2796], RIGHT_GRAPH[2732], RIGHT_GRAPH[2668], RIGHT_GRAPH[2604]};
					9'd365	:	PATTERN = {RIGHT_GRAPH[3053], RIGHT_GRAPH[2989], RIGHT_GRAPH[2925], RIGHT_GRAPH[2861], RIGHT_GRAPH[2797], RIGHT_GRAPH[2733], RIGHT_GRAPH[2669], RIGHT_GRAPH[2605]};
					9'd366	:	PATTERN = {RIGHT_GRAPH[3054], RIGHT_GRAPH[2990], RIGHT_GRAPH[2926], RIGHT_GRAPH[2862], RIGHT_GRAPH[2798], RIGHT_GRAPH[2734], RIGHT_GRAPH[2670], RIGHT_GRAPH[2606]};
					9'd367	:	PATTERN = {RIGHT_GRAPH[3055], RIGHT_GRAPH[2991], RIGHT_GRAPH[2927], RIGHT_GRAPH[2863], RIGHT_GRAPH[2799], RIGHT_GRAPH[2735], RIGHT_GRAPH[2671], RIGHT_GRAPH[2607]};
					9'd368	:	PATTERN = {RIGHT_GRAPH[3056], RIGHT_GRAPH[2992], RIGHT_GRAPH[2928], RIGHT_GRAPH[2864], RIGHT_GRAPH[2800], RIGHT_GRAPH[2736], RIGHT_GRAPH[2672], RIGHT_GRAPH[2608]};
					9'd369	:	PATTERN = {RIGHT_GRAPH[3057], RIGHT_GRAPH[2993], RIGHT_GRAPH[2929], RIGHT_GRAPH[2865], RIGHT_GRAPH[2801], RIGHT_GRAPH[2737], RIGHT_GRAPH[2673], RIGHT_GRAPH[2609]};
					9'd370	:	PATTERN = {RIGHT_GRAPH[3058], RIGHT_GRAPH[2994], RIGHT_GRAPH[2930], RIGHT_GRAPH[2866], RIGHT_GRAPH[2802], RIGHT_GRAPH[2738], RIGHT_GRAPH[2674], RIGHT_GRAPH[2610]};
					9'd371	:	PATTERN = {RIGHT_GRAPH[3059], RIGHT_GRAPH[2995], RIGHT_GRAPH[2931], RIGHT_GRAPH[2867], RIGHT_GRAPH[2803], RIGHT_GRAPH[2739], RIGHT_GRAPH[2675], RIGHT_GRAPH[2611]};
					9'd372	:	PATTERN = {RIGHT_GRAPH[3060], RIGHT_GRAPH[2996], RIGHT_GRAPH[2932], RIGHT_GRAPH[2868], RIGHT_GRAPH[2804], RIGHT_GRAPH[2740], RIGHT_GRAPH[2676], RIGHT_GRAPH[2612]};
					9'd373	:	PATTERN = {RIGHT_GRAPH[3061], RIGHT_GRAPH[2997], RIGHT_GRAPH[2933], RIGHT_GRAPH[2869], RIGHT_GRAPH[2805], RIGHT_GRAPH[2741], RIGHT_GRAPH[2677], RIGHT_GRAPH[2613]};
					9'd374	:	PATTERN = {RIGHT_GRAPH[3062], RIGHT_GRAPH[2998], RIGHT_GRAPH[2934], RIGHT_GRAPH[2870], RIGHT_GRAPH[2806], RIGHT_GRAPH[2742], RIGHT_GRAPH[2678], RIGHT_GRAPH[2614]};
					9'd375	:	PATTERN = {RIGHT_GRAPH[3063], RIGHT_GRAPH[2999], RIGHT_GRAPH[2935], RIGHT_GRAPH[2871], RIGHT_GRAPH[2807], RIGHT_GRAPH[2743], RIGHT_GRAPH[2679], RIGHT_GRAPH[2615]};
					9'd376	:	PATTERN = {RIGHT_GRAPH[3064], RIGHT_GRAPH[3000], RIGHT_GRAPH[2936], RIGHT_GRAPH[2872], RIGHT_GRAPH[2808], RIGHT_GRAPH[2744], RIGHT_GRAPH[2680], RIGHT_GRAPH[2616]};
					9'd377	:	PATTERN = {RIGHT_GRAPH[3065], RIGHT_GRAPH[3001], RIGHT_GRAPH[2937], RIGHT_GRAPH[2873], RIGHT_GRAPH[2809], RIGHT_GRAPH[2745], RIGHT_GRAPH[2681], RIGHT_GRAPH[2617]};
					9'd378	:	PATTERN = {RIGHT_GRAPH[3066], RIGHT_GRAPH[3002], RIGHT_GRAPH[2938], RIGHT_GRAPH[2874], RIGHT_GRAPH[2810], RIGHT_GRAPH[2746], RIGHT_GRAPH[2682], RIGHT_GRAPH[2618]};
					9'd379	:	PATTERN = {RIGHT_GRAPH[3067], RIGHT_GRAPH[3003], RIGHT_GRAPH[2939], RIGHT_GRAPH[2875], RIGHT_GRAPH[2811], RIGHT_GRAPH[2747], RIGHT_GRAPH[2683], RIGHT_GRAPH[2619]};
					9'd380	:	PATTERN = {RIGHT_GRAPH[3068], RIGHT_GRAPH[3004], RIGHT_GRAPH[2940], RIGHT_GRAPH[2876], RIGHT_GRAPH[2812], RIGHT_GRAPH[2748], RIGHT_GRAPH[2684], RIGHT_GRAPH[2620]};
					9'd381	:	PATTERN = {RIGHT_GRAPH[3069], RIGHT_GRAPH[3005], RIGHT_GRAPH[2941], RIGHT_GRAPH[2877], RIGHT_GRAPH[2813], RIGHT_GRAPH[2749], RIGHT_GRAPH[2685], RIGHT_GRAPH[2621]};
					9'd382	:	PATTERN = {RIGHT_GRAPH[3070], RIGHT_GRAPH[3006], RIGHT_GRAPH[2942], RIGHT_GRAPH[2878], RIGHT_GRAPH[2814], RIGHT_GRAPH[2750], RIGHT_GRAPH[2686], RIGHT_GRAPH[2622]};
					9'd383	:	PATTERN = {RIGHT_GRAPH[3071], RIGHT_GRAPH[3007], RIGHT_GRAPH[2943], RIGHT_GRAPH[2879], RIGHT_GRAPH[2815], RIGHT_GRAPH[2751], RIGHT_GRAPH[2687], RIGHT_GRAPH[2623]};
					9'd384	:	PATTERN = {RIGHT_GRAPH[3520], RIGHT_GRAPH[3456], RIGHT_GRAPH[3392], RIGHT_GRAPH[3328], RIGHT_GRAPH[3264], RIGHT_GRAPH[3200], RIGHT_GRAPH[3136], RIGHT_GRAPH[3072]};
					9'd385	:	PATTERN = {RIGHT_GRAPH[3521], RIGHT_GRAPH[3457], RIGHT_GRAPH[3393], RIGHT_GRAPH[3329], RIGHT_GRAPH[3265], RIGHT_GRAPH[3201], RIGHT_GRAPH[3137], RIGHT_GRAPH[3073]};
					9'd386	:	PATTERN = {RIGHT_GRAPH[3522], RIGHT_GRAPH[3458], RIGHT_GRAPH[3394], RIGHT_GRAPH[3330], RIGHT_GRAPH[3266], RIGHT_GRAPH[3202], RIGHT_GRAPH[3138], RIGHT_GRAPH[3074]};
					9'd387	:	PATTERN = {RIGHT_GRAPH[3523], RIGHT_GRAPH[3459], RIGHT_GRAPH[3395], RIGHT_GRAPH[3331], RIGHT_GRAPH[3267], RIGHT_GRAPH[3203], RIGHT_GRAPH[3139], RIGHT_GRAPH[3075]};
					9'd388	:	PATTERN = {RIGHT_GRAPH[3524], RIGHT_GRAPH[3460], RIGHT_GRAPH[3396], RIGHT_GRAPH[3332], RIGHT_GRAPH[3268], RIGHT_GRAPH[3204], RIGHT_GRAPH[3140], RIGHT_GRAPH[3076]};
					9'd389	:	PATTERN = {RIGHT_GRAPH[3525], RIGHT_GRAPH[3461], RIGHT_GRAPH[3397], RIGHT_GRAPH[3333], RIGHT_GRAPH[3269], RIGHT_GRAPH[3205], RIGHT_GRAPH[3141], RIGHT_GRAPH[3077]};
					9'd390	:	PATTERN = {RIGHT_GRAPH[3526], RIGHT_GRAPH[3462], RIGHT_GRAPH[3398], RIGHT_GRAPH[3334], RIGHT_GRAPH[3270], RIGHT_GRAPH[3206], RIGHT_GRAPH[3142], RIGHT_GRAPH[3078]};
					9'd391	:	PATTERN = {RIGHT_GRAPH[3527], RIGHT_GRAPH[3463], RIGHT_GRAPH[3399], RIGHT_GRAPH[3335], RIGHT_GRAPH[3271], RIGHT_GRAPH[3207], RIGHT_GRAPH[3143], RIGHT_GRAPH[3079]};
					9'd392	:	PATTERN = {RIGHT_GRAPH[3528], RIGHT_GRAPH[3464], RIGHT_GRAPH[3400], RIGHT_GRAPH[3336], RIGHT_GRAPH[3272], RIGHT_GRAPH[3208], RIGHT_GRAPH[3144], RIGHT_GRAPH[3080]};
					9'd393	:	PATTERN = {RIGHT_GRAPH[3529], RIGHT_GRAPH[3465], RIGHT_GRAPH[3401], RIGHT_GRAPH[3337], RIGHT_GRAPH[3273], RIGHT_GRAPH[3209], RIGHT_GRAPH[3145], RIGHT_GRAPH[3081]};
					9'd394	:	PATTERN = {RIGHT_GRAPH[3530], RIGHT_GRAPH[3466], RIGHT_GRAPH[3402], RIGHT_GRAPH[3338], RIGHT_GRAPH[3274], RIGHT_GRAPH[3210], RIGHT_GRAPH[3146], RIGHT_GRAPH[3082]};
					9'd395	:	PATTERN = {RIGHT_GRAPH[3531], RIGHT_GRAPH[3467], RIGHT_GRAPH[3403], RIGHT_GRAPH[3339], RIGHT_GRAPH[3275], RIGHT_GRAPH[3211], RIGHT_GRAPH[3147], RIGHT_GRAPH[3083]};
					9'd396	:	PATTERN = {RIGHT_GRAPH[3532], RIGHT_GRAPH[3468], RIGHT_GRAPH[3404], RIGHT_GRAPH[3340], RIGHT_GRAPH[3276], RIGHT_GRAPH[3212], RIGHT_GRAPH[3148], RIGHT_GRAPH[3084]};
					9'd397	:	PATTERN = {RIGHT_GRAPH[3533], RIGHT_GRAPH[3469], RIGHT_GRAPH[3405], RIGHT_GRAPH[3341], RIGHT_GRAPH[3277], RIGHT_GRAPH[3213], RIGHT_GRAPH[3149], RIGHT_GRAPH[3085]};
					9'd398	:	PATTERN = {RIGHT_GRAPH[3534], RIGHT_GRAPH[3470], RIGHT_GRAPH[3406], RIGHT_GRAPH[3342], RIGHT_GRAPH[3278], RIGHT_GRAPH[3214], RIGHT_GRAPH[3150], RIGHT_GRAPH[3086]};
					9'd399	:	PATTERN = {RIGHT_GRAPH[3535], RIGHT_GRAPH[3471], RIGHT_GRAPH[3407], RIGHT_GRAPH[3343], RIGHT_GRAPH[3279], RIGHT_GRAPH[3215], RIGHT_GRAPH[3151], RIGHT_GRAPH[3087]};
					9'd400	:	PATTERN = {RIGHT_GRAPH[3536], RIGHT_GRAPH[3472], RIGHT_GRAPH[3408], RIGHT_GRAPH[3344], RIGHT_GRAPH[3280], RIGHT_GRAPH[3216], RIGHT_GRAPH[3152], RIGHT_GRAPH[3088]};
					9'd401	:	PATTERN = {RIGHT_GRAPH[3537], RIGHT_GRAPH[3473], RIGHT_GRAPH[3409], RIGHT_GRAPH[3345], RIGHT_GRAPH[3281], RIGHT_GRAPH[3217], RIGHT_GRAPH[3153], RIGHT_GRAPH[3089]};
					9'd402	:	PATTERN = {RIGHT_GRAPH[3538], RIGHT_GRAPH[3474], RIGHT_GRAPH[3410], RIGHT_GRAPH[3346], RIGHT_GRAPH[3282], RIGHT_GRAPH[3218], RIGHT_GRAPH[3154], RIGHT_GRAPH[3090]};
					9'd403	:	PATTERN = {RIGHT_GRAPH[3539], RIGHT_GRAPH[3475], RIGHT_GRAPH[3411], RIGHT_GRAPH[3347], RIGHT_GRAPH[3283], RIGHT_GRAPH[3219], RIGHT_GRAPH[3155], RIGHT_GRAPH[3091]};
					9'd404	:	PATTERN = {RIGHT_GRAPH[3540], RIGHT_GRAPH[3476], RIGHT_GRAPH[3412], RIGHT_GRAPH[3348], RIGHT_GRAPH[3284], RIGHT_GRAPH[3220], RIGHT_GRAPH[3156], RIGHT_GRAPH[3092]};
					9'd405	:	PATTERN = {RIGHT_GRAPH[3541], RIGHT_GRAPH[3477], RIGHT_GRAPH[3413], RIGHT_GRAPH[3349], RIGHT_GRAPH[3285], RIGHT_GRAPH[3221], RIGHT_GRAPH[3157], RIGHT_GRAPH[3093]};
					9'd406	:	PATTERN = {RIGHT_GRAPH[3542], RIGHT_GRAPH[3478], RIGHT_GRAPH[3414], RIGHT_GRAPH[3350], RIGHT_GRAPH[3286], RIGHT_GRAPH[3222], RIGHT_GRAPH[3158], RIGHT_GRAPH[3094]};
					9'd407	:	PATTERN = {RIGHT_GRAPH[3543], RIGHT_GRAPH[3479], RIGHT_GRAPH[3415], RIGHT_GRAPH[3351], RIGHT_GRAPH[3287], RIGHT_GRAPH[3223], RIGHT_GRAPH[3159], RIGHT_GRAPH[3095]};
					9'd408	:	PATTERN = {RIGHT_GRAPH[3544], RIGHT_GRAPH[3480], RIGHT_GRAPH[3416], RIGHT_GRAPH[3352], RIGHT_GRAPH[3288], RIGHT_GRAPH[3224], RIGHT_GRAPH[3160], RIGHT_GRAPH[3096]};
					9'd409	:	PATTERN = {RIGHT_GRAPH[3545], RIGHT_GRAPH[3481], RIGHT_GRAPH[3417], RIGHT_GRAPH[3353], RIGHT_GRAPH[3289], RIGHT_GRAPH[3225], RIGHT_GRAPH[3161], RIGHT_GRAPH[3097]};
					9'd410	:	PATTERN = {RIGHT_GRAPH[3546], RIGHT_GRAPH[3482], RIGHT_GRAPH[3418], RIGHT_GRAPH[3354], RIGHT_GRAPH[3290], RIGHT_GRAPH[3226], RIGHT_GRAPH[3162], RIGHT_GRAPH[3098]};
					9'd411	:	PATTERN = {RIGHT_GRAPH[3547], RIGHT_GRAPH[3483], RIGHT_GRAPH[3419], RIGHT_GRAPH[3355], RIGHT_GRAPH[3291], RIGHT_GRAPH[3227], RIGHT_GRAPH[3163], RIGHT_GRAPH[3099]};
					9'd412	:	PATTERN = {RIGHT_GRAPH[3548], RIGHT_GRAPH[3484], RIGHT_GRAPH[3420], RIGHT_GRAPH[3356], RIGHT_GRAPH[3292], RIGHT_GRAPH[3228], RIGHT_GRAPH[3164], RIGHT_GRAPH[3100]};
					9'd413	:	PATTERN = {RIGHT_GRAPH[3549], RIGHT_GRAPH[3485], RIGHT_GRAPH[3421], RIGHT_GRAPH[3357], RIGHT_GRAPH[3293], RIGHT_GRAPH[3229], RIGHT_GRAPH[3165], RIGHT_GRAPH[3101]};
					9'd414	:	PATTERN = {RIGHT_GRAPH[3550], RIGHT_GRAPH[3486], RIGHT_GRAPH[3422], RIGHT_GRAPH[3358], RIGHT_GRAPH[3294], RIGHT_GRAPH[3230], RIGHT_GRAPH[3166], RIGHT_GRAPH[3102]};
					9'd415	:	PATTERN = {RIGHT_GRAPH[3551], RIGHT_GRAPH[3487], RIGHT_GRAPH[3423], RIGHT_GRAPH[3359], RIGHT_GRAPH[3295], RIGHT_GRAPH[3231], RIGHT_GRAPH[3167], RIGHT_GRAPH[3103]};
					9'd416	:	PATTERN = {RIGHT_GRAPH[3552], RIGHT_GRAPH[3488], RIGHT_GRAPH[3424], RIGHT_GRAPH[3360], RIGHT_GRAPH[3296], RIGHT_GRAPH[3232], RIGHT_GRAPH[3168], RIGHT_GRAPH[3104]};
					9'd417	:	PATTERN = {RIGHT_GRAPH[3553], RIGHT_GRAPH[3489], RIGHT_GRAPH[3425], RIGHT_GRAPH[3361], RIGHT_GRAPH[3297], RIGHT_GRAPH[3233], RIGHT_GRAPH[3169], RIGHT_GRAPH[3105]};
					9'd418	:	PATTERN = {RIGHT_GRAPH[3554], RIGHT_GRAPH[3490], RIGHT_GRAPH[3426], RIGHT_GRAPH[3362], RIGHT_GRAPH[3298], RIGHT_GRAPH[3234], RIGHT_GRAPH[3170], RIGHT_GRAPH[3106]};
					9'd419	:	PATTERN = {RIGHT_GRAPH[3555], RIGHT_GRAPH[3491], RIGHT_GRAPH[3427], RIGHT_GRAPH[3363], RIGHT_GRAPH[3299], RIGHT_GRAPH[3235], RIGHT_GRAPH[3171], RIGHT_GRAPH[3107]};
					9'd420	:	PATTERN = {RIGHT_GRAPH[3556], RIGHT_GRAPH[3492], RIGHT_GRAPH[3428], RIGHT_GRAPH[3364], RIGHT_GRAPH[3300], RIGHT_GRAPH[3236], RIGHT_GRAPH[3172], RIGHT_GRAPH[3108]};
					9'd421	:	PATTERN = {RIGHT_GRAPH[3557], RIGHT_GRAPH[3493], RIGHT_GRAPH[3429], RIGHT_GRAPH[3365], RIGHT_GRAPH[3301], RIGHT_GRAPH[3237], RIGHT_GRAPH[3173], RIGHT_GRAPH[3109]};
					9'd422	:	PATTERN = {RIGHT_GRAPH[3558], RIGHT_GRAPH[3494], RIGHT_GRAPH[3430], RIGHT_GRAPH[3366], RIGHT_GRAPH[3302], RIGHT_GRAPH[3238], RIGHT_GRAPH[3174], RIGHT_GRAPH[3110]};
					9'd423	:	PATTERN = {RIGHT_GRAPH[3559], RIGHT_GRAPH[3495], RIGHT_GRAPH[3431], RIGHT_GRAPH[3367], RIGHT_GRAPH[3303], RIGHT_GRAPH[3239], RIGHT_GRAPH[3175], RIGHT_GRAPH[3111]};
					9'd424	:	PATTERN = {RIGHT_GRAPH[3560], RIGHT_GRAPH[3496], RIGHT_GRAPH[3432], RIGHT_GRAPH[3368], RIGHT_GRAPH[3304], RIGHT_GRAPH[3240], RIGHT_GRAPH[3176], RIGHT_GRAPH[3112]};
					9'd425	:	PATTERN = {RIGHT_GRAPH[3561], RIGHT_GRAPH[3497], RIGHT_GRAPH[3433], RIGHT_GRAPH[3369], RIGHT_GRAPH[3305], RIGHT_GRAPH[3241], RIGHT_GRAPH[3177], RIGHT_GRAPH[3113]};
					9'd426	:	PATTERN = {RIGHT_GRAPH[3562], RIGHT_GRAPH[3498], RIGHT_GRAPH[3434], RIGHT_GRAPH[3370], RIGHT_GRAPH[3306], RIGHT_GRAPH[3242], RIGHT_GRAPH[3178], RIGHT_GRAPH[3114]};
					9'd427	:	PATTERN = {RIGHT_GRAPH[3563], RIGHT_GRAPH[3499], RIGHT_GRAPH[3435], RIGHT_GRAPH[3371], RIGHT_GRAPH[3307], RIGHT_GRAPH[3243], RIGHT_GRAPH[3179], RIGHT_GRAPH[3115]};
					9'd428	:	PATTERN = {RIGHT_GRAPH[3564], RIGHT_GRAPH[3500], RIGHT_GRAPH[3436], RIGHT_GRAPH[3372], RIGHT_GRAPH[3308], RIGHT_GRAPH[3244], RIGHT_GRAPH[3180], RIGHT_GRAPH[3116]};
					9'd429	:	PATTERN = {RIGHT_GRAPH[3565], RIGHT_GRAPH[3501], RIGHT_GRAPH[3437], RIGHT_GRAPH[3373], RIGHT_GRAPH[3309], RIGHT_GRAPH[3245], RIGHT_GRAPH[3181], RIGHT_GRAPH[3117]};
					9'd430	:	PATTERN = {RIGHT_GRAPH[3566], RIGHT_GRAPH[3502], RIGHT_GRAPH[3438], RIGHT_GRAPH[3374], RIGHT_GRAPH[3310], RIGHT_GRAPH[3246], RIGHT_GRAPH[3182], RIGHT_GRAPH[3118]};
					9'd431	:	PATTERN = {RIGHT_GRAPH[3567], RIGHT_GRAPH[3503], RIGHT_GRAPH[3439], RIGHT_GRAPH[3375], RIGHT_GRAPH[3311], RIGHT_GRAPH[3247], RIGHT_GRAPH[3183], RIGHT_GRAPH[3119]};
					9'd432	:	PATTERN = {RIGHT_GRAPH[3568], RIGHT_GRAPH[3504], RIGHT_GRAPH[3440], RIGHT_GRAPH[3376], RIGHT_GRAPH[3312], RIGHT_GRAPH[3248], RIGHT_GRAPH[3184], RIGHT_GRAPH[3120]};
					9'd433	:	PATTERN = {RIGHT_GRAPH[3569], RIGHT_GRAPH[3505], RIGHT_GRAPH[3441], RIGHT_GRAPH[3377], RIGHT_GRAPH[3313], RIGHT_GRAPH[3249], RIGHT_GRAPH[3185], RIGHT_GRAPH[3121]};
					9'd434	:	PATTERN = {RIGHT_GRAPH[3570], RIGHT_GRAPH[3506], RIGHT_GRAPH[3442], RIGHT_GRAPH[3378], RIGHT_GRAPH[3314], RIGHT_GRAPH[3250], RIGHT_GRAPH[3186], RIGHT_GRAPH[3122]};
					9'd435	:	PATTERN = {RIGHT_GRAPH[3571], RIGHT_GRAPH[3507], RIGHT_GRAPH[3443], RIGHT_GRAPH[3379], RIGHT_GRAPH[3315], RIGHT_GRAPH[3251], RIGHT_GRAPH[3187], RIGHT_GRAPH[3123]};
					9'd436	:	PATTERN = {RIGHT_GRAPH[3572], RIGHT_GRAPH[3508], RIGHT_GRAPH[3444], RIGHT_GRAPH[3380], RIGHT_GRAPH[3316], RIGHT_GRAPH[3252], RIGHT_GRAPH[3188], RIGHT_GRAPH[3124]};
					9'd437	:	PATTERN = {RIGHT_GRAPH[3573], RIGHT_GRAPH[3509], RIGHT_GRAPH[3445], RIGHT_GRAPH[3381], RIGHT_GRAPH[3317], RIGHT_GRAPH[3253], RIGHT_GRAPH[3189], RIGHT_GRAPH[3125]};
					9'd438	:	PATTERN = {RIGHT_GRAPH[3574], RIGHT_GRAPH[3510], RIGHT_GRAPH[3446], RIGHT_GRAPH[3382], RIGHT_GRAPH[3318], RIGHT_GRAPH[3254], RIGHT_GRAPH[3190], RIGHT_GRAPH[3126]};
					9'd439	:	PATTERN = {RIGHT_GRAPH[3575], RIGHT_GRAPH[3511], RIGHT_GRAPH[3447], RIGHT_GRAPH[3383], RIGHT_GRAPH[3319], RIGHT_GRAPH[3255], RIGHT_GRAPH[3191], RIGHT_GRAPH[3127]};
					9'd440	:	PATTERN = {RIGHT_GRAPH[3576], RIGHT_GRAPH[3512], RIGHT_GRAPH[3448], RIGHT_GRAPH[3384], RIGHT_GRAPH[3320], RIGHT_GRAPH[3256], RIGHT_GRAPH[3192], RIGHT_GRAPH[3128]};
					9'd441	:	PATTERN = {RIGHT_GRAPH[3577], RIGHT_GRAPH[3513], RIGHT_GRAPH[3449], RIGHT_GRAPH[3385], RIGHT_GRAPH[3321], RIGHT_GRAPH[3257], RIGHT_GRAPH[3193], RIGHT_GRAPH[3129]};
					9'd442	:	PATTERN = {RIGHT_GRAPH[3578], RIGHT_GRAPH[3514], RIGHT_GRAPH[3450], RIGHT_GRAPH[3386], RIGHT_GRAPH[3322], RIGHT_GRAPH[3258], RIGHT_GRAPH[3194], RIGHT_GRAPH[3130]};
					9'd443	:	PATTERN = {RIGHT_GRAPH[3579], RIGHT_GRAPH[3515], RIGHT_GRAPH[3451], RIGHT_GRAPH[3387], RIGHT_GRAPH[3323], RIGHT_GRAPH[3259], RIGHT_GRAPH[3195], RIGHT_GRAPH[3131]};
					9'd444	:	PATTERN = {RIGHT_GRAPH[3580], RIGHT_GRAPH[3516], RIGHT_GRAPH[3452], RIGHT_GRAPH[3388], RIGHT_GRAPH[3324], RIGHT_GRAPH[3260], RIGHT_GRAPH[3196], RIGHT_GRAPH[3132]};
					9'd445	:	PATTERN = {RIGHT_GRAPH[3581], RIGHT_GRAPH[3517], RIGHT_GRAPH[3453], RIGHT_GRAPH[3389], RIGHT_GRAPH[3325], RIGHT_GRAPH[3261], RIGHT_GRAPH[3197], RIGHT_GRAPH[3133]};
					9'd446	:	PATTERN = {RIGHT_GRAPH[3582], RIGHT_GRAPH[3518], RIGHT_GRAPH[3454], RIGHT_GRAPH[3390], RIGHT_GRAPH[3326], RIGHT_GRAPH[3262], RIGHT_GRAPH[3198], RIGHT_GRAPH[3134]};
					9'd447	:	PATTERN = {RIGHT_GRAPH[3583], RIGHT_GRAPH[3519], RIGHT_GRAPH[3455], RIGHT_GRAPH[3391], RIGHT_GRAPH[3327], RIGHT_GRAPH[3263], RIGHT_GRAPH[3199], RIGHT_GRAPH[3135]};
					9'd448	:	PATTERN = {RIGHT_GRAPH[4032], RIGHT_GRAPH[3968], RIGHT_GRAPH[3904], RIGHT_GRAPH[3840], RIGHT_GRAPH[3776], RIGHT_GRAPH[3712], RIGHT_GRAPH[3648], RIGHT_GRAPH[3584]};
					9'd449	:	PATTERN = {RIGHT_GRAPH[4033], RIGHT_GRAPH[3969], RIGHT_GRAPH[3905], RIGHT_GRAPH[3841], RIGHT_GRAPH[3777], RIGHT_GRAPH[3713], RIGHT_GRAPH[3649], RIGHT_GRAPH[3585]};
					9'd450	:	PATTERN = {RIGHT_GRAPH[4034], RIGHT_GRAPH[3970], RIGHT_GRAPH[3906], RIGHT_GRAPH[3842], RIGHT_GRAPH[3778], RIGHT_GRAPH[3714], RIGHT_GRAPH[3650], RIGHT_GRAPH[3586]};
					9'd451	:	PATTERN = {RIGHT_GRAPH[4035], RIGHT_GRAPH[3971], RIGHT_GRAPH[3907], RIGHT_GRAPH[3843], RIGHT_GRAPH[3779], RIGHT_GRAPH[3715], RIGHT_GRAPH[3651], RIGHT_GRAPH[3587]};
					9'd452	:	PATTERN = {RIGHT_GRAPH[4036], RIGHT_GRAPH[3972], RIGHT_GRAPH[3908], RIGHT_GRAPH[3844], RIGHT_GRAPH[3780], RIGHT_GRAPH[3716], RIGHT_GRAPH[3652], RIGHT_GRAPH[3588]};
					9'd453	:	PATTERN = {RIGHT_GRAPH[4037], RIGHT_GRAPH[3973], RIGHT_GRAPH[3909], RIGHT_GRAPH[3845], RIGHT_GRAPH[3781], RIGHT_GRAPH[3717], RIGHT_GRAPH[3653], RIGHT_GRAPH[3589]};
					9'd454	:	PATTERN = {RIGHT_GRAPH[4038], RIGHT_GRAPH[3974], RIGHT_GRAPH[3910], RIGHT_GRAPH[3846], RIGHT_GRAPH[3782], RIGHT_GRAPH[3718], RIGHT_GRAPH[3654], RIGHT_GRAPH[3590]};
					9'd455	:	PATTERN = {RIGHT_GRAPH[4039], RIGHT_GRAPH[3975], RIGHT_GRAPH[3911], RIGHT_GRAPH[3847], RIGHT_GRAPH[3783], RIGHT_GRAPH[3719], RIGHT_GRAPH[3655], RIGHT_GRAPH[3591]};
					9'd456	:	PATTERN = {RIGHT_GRAPH[4040], RIGHT_GRAPH[3976], RIGHT_GRAPH[3912], RIGHT_GRAPH[3848], RIGHT_GRAPH[3784], RIGHT_GRAPH[3720], RIGHT_GRAPH[3656], RIGHT_GRAPH[3592]};
					9'd457	:	PATTERN = {RIGHT_GRAPH[4041], RIGHT_GRAPH[3977], RIGHT_GRAPH[3913], RIGHT_GRAPH[3849], RIGHT_GRAPH[3785], RIGHT_GRAPH[3721], RIGHT_GRAPH[3657], RIGHT_GRAPH[3593]};
					9'd458	:	PATTERN = {RIGHT_GRAPH[4042], RIGHT_GRAPH[3978], RIGHT_GRAPH[3914], RIGHT_GRAPH[3850], RIGHT_GRAPH[3786], RIGHT_GRAPH[3722], RIGHT_GRAPH[3658], RIGHT_GRAPH[3594]};
					9'd459	:	PATTERN = {RIGHT_GRAPH[4043], RIGHT_GRAPH[3979], RIGHT_GRAPH[3915], RIGHT_GRAPH[3851], RIGHT_GRAPH[3787], RIGHT_GRAPH[3723], RIGHT_GRAPH[3659], RIGHT_GRAPH[3595]};
					9'd460	:	PATTERN = {RIGHT_GRAPH[4044], RIGHT_GRAPH[3980], RIGHT_GRAPH[3916], RIGHT_GRAPH[3852], RIGHT_GRAPH[3788], RIGHT_GRAPH[3724], RIGHT_GRAPH[3660], RIGHT_GRAPH[3596]};
					9'd461	:	PATTERN = {RIGHT_GRAPH[4045], RIGHT_GRAPH[3981], RIGHT_GRAPH[3917], RIGHT_GRAPH[3853], RIGHT_GRAPH[3789], RIGHT_GRAPH[3725], RIGHT_GRAPH[3661], RIGHT_GRAPH[3597]};
					9'd462	:	PATTERN = {RIGHT_GRAPH[4046], RIGHT_GRAPH[3982], RIGHT_GRAPH[3918], RIGHT_GRAPH[3854], RIGHT_GRAPH[3790], RIGHT_GRAPH[3726], RIGHT_GRAPH[3662], RIGHT_GRAPH[3598]};
					9'd463	:	PATTERN = {RIGHT_GRAPH[4047], RIGHT_GRAPH[3983], RIGHT_GRAPH[3919], RIGHT_GRAPH[3855], RIGHT_GRAPH[3791], RIGHT_GRAPH[3727], RIGHT_GRAPH[3663], RIGHT_GRAPH[3599]};
					9'd464	:	PATTERN = {RIGHT_GRAPH[4048], RIGHT_GRAPH[3984], RIGHT_GRAPH[3920], RIGHT_GRAPH[3856], RIGHT_GRAPH[3792], RIGHT_GRAPH[3728], RIGHT_GRAPH[3664], RIGHT_GRAPH[3600]};
					9'd465	:	PATTERN = {RIGHT_GRAPH[4049], RIGHT_GRAPH[3985], RIGHT_GRAPH[3921], RIGHT_GRAPH[3857], RIGHT_GRAPH[3793], RIGHT_GRAPH[3729], RIGHT_GRAPH[3665], RIGHT_GRAPH[3601]};
					9'd466	:	PATTERN = {RIGHT_GRAPH[4050], RIGHT_GRAPH[3986], RIGHT_GRAPH[3922], RIGHT_GRAPH[3858], RIGHT_GRAPH[3794], RIGHT_GRAPH[3730], RIGHT_GRAPH[3666], RIGHT_GRAPH[3602]};
					9'd467	:	PATTERN = {RIGHT_GRAPH[4051], RIGHT_GRAPH[3987], RIGHT_GRAPH[3923], RIGHT_GRAPH[3859], RIGHT_GRAPH[3795], RIGHT_GRAPH[3731], RIGHT_GRAPH[3667], RIGHT_GRAPH[3603]};
					9'd468	:	PATTERN = {RIGHT_GRAPH[4052], RIGHT_GRAPH[3988], RIGHT_GRAPH[3924], RIGHT_GRAPH[3860], RIGHT_GRAPH[3796], RIGHT_GRAPH[3732], RIGHT_GRAPH[3668], RIGHT_GRAPH[3604]};
					9'd469	:	PATTERN = {RIGHT_GRAPH[4053], RIGHT_GRAPH[3989], RIGHT_GRAPH[3925], RIGHT_GRAPH[3861], RIGHT_GRAPH[3797], RIGHT_GRAPH[3733], RIGHT_GRAPH[3669], RIGHT_GRAPH[3605]};
					9'd470	:	PATTERN = {RIGHT_GRAPH[4054], RIGHT_GRAPH[3990], RIGHT_GRAPH[3926], RIGHT_GRAPH[3862], RIGHT_GRAPH[3798], RIGHT_GRAPH[3734], RIGHT_GRAPH[3670], RIGHT_GRAPH[3606]};
					9'd471	:	PATTERN = {RIGHT_GRAPH[4055], RIGHT_GRAPH[3991], RIGHT_GRAPH[3927], RIGHT_GRAPH[3863], RIGHT_GRAPH[3799], RIGHT_GRAPH[3735], RIGHT_GRAPH[3671], RIGHT_GRAPH[3607]};
					9'd472	:	PATTERN = {RIGHT_GRAPH[4056], RIGHT_GRAPH[3992], RIGHT_GRAPH[3928], RIGHT_GRAPH[3864], RIGHT_GRAPH[3800], RIGHT_GRAPH[3736], RIGHT_GRAPH[3672], RIGHT_GRAPH[3608]};
					9'd473	:	PATTERN = {RIGHT_GRAPH[4057], RIGHT_GRAPH[3993], RIGHT_GRAPH[3929], RIGHT_GRAPH[3865], RIGHT_GRAPH[3801], RIGHT_GRAPH[3737], RIGHT_GRAPH[3673], RIGHT_GRAPH[3609]};
					9'd474	:	PATTERN = {RIGHT_GRAPH[4058], RIGHT_GRAPH[3994], RIGHT_GRAPH[3930], RIGHT_GRAPH[3866], RIGHT_GRAPH[3802], RIGHT_GRAPH[3738], RIGHT_GRAPH[3674], RIGHT_GRAPH[3610]};
					9'd475	:	PATTERN = {RIGHT_GRAPH[4059], RIGHT_GRAPH[3995], RIGHT_GRAPH[3931], RIGHT_GRAPH[3867], RIGHT_GRAPH[3803], RIGHT_GRAPH[3739], RIGHT_GRAPH[3675], RIGHT_GRAPH[3611]};
					9'd476	:	PATTERN = {RIGHT_GRAPH[4060], RIGHT_GRAPH[3996], RIGHT_GRAPH[3932], RIGHT_GRAPH[3868], RIGHT_GRAPH[3804], RIGHT_GRAPH[3740], RIGHT_GRAPH[3676], RIGHT_GRAPH[3612]};
					9'd477	:	PATTERN = {RIGHT_GRAPH[4061], RIGHT_GRAPH[3997], RIGHT_GRAPH[3933], RIGHT_GRAPH[3869], RIGHT_GRAPH[3805], RIGHT_GRAPH[3741], RIGHT_GRAPH[3677], RIGHT_GRAPH[3613]};
					9'd478	:	PATTERN = {RIGHT_GRAPH[4062], RIGHT_GRAPH[3998], RIGHT_GRAPH[3934], RIGHT_GRAPH[3870], RIGHT_GRAPH[3806], RIGHT_GRAPH[3742], RIGHT_GRAPH[3678], RIGHT_GRAPH[3614]};
					9'd479	:	PATTERN = {RIGHT_GRAPH[4063], RIGHT_GRAPH[3999], RIGHT_GRAPH[3935], RIGHT_GRAPH[3871], RIGHT_GRAPH[3807], RIGHT_GRAPH[3743], RIGHT_GRAPH[3679], RIGHT_GRAPH[3615]};
					9'd480	:	PATTERN = {RIGHT_GRAPH[4064], RIGHT_GRAPH[4000], RIGHT_GRAPH[3936], RIGHT_GRAPH[3872], RIGHT_GRAPH[3808], RIGHT_GRAPH[3744], RIGHT_GRAPH[3680], RIGHT_GRAPH[3616]};
					9'd481	:	PATTERN = {RIGHT_GRAPH[4065], RIGHT_GRAPH[4001], RIGHT_GRAPH[3937], RIGHT_GRAPH[3873], RIGHT_GRAPH[3809], RIGHT_GRAPH[3745], RIGHT_GRAPH[3681], RIGHT_GRAPH[3617]};
					9'd482	:	PATTERN = {RIGHT_GRAPH[4066], RIGHT_GRAPH[4002], RIGHT_GRAPH[3938], RIGHT_GRAPH[3874], RIGHT_GRAPH[3810], RIGHT_GRAPH[3746], RIGHT_GRAPH[3682], RIGHT_GRAPH[3618]};
					9'd483	:	PATTERN = {RIGHT_GRAPH[4067], RIGHT_GRAPH[4003], RIGHT_GRAPH[3939], RIGHT_GRAPH[3875], RIGHT_GRAPH[3811], RIGHT_GRAPH[3747], RIGHT_GRAPH[3683], RIGHT_GRAPH[3619]};
					9'd484	:	PATTERN = {RIGHT_GRAPH[4068], RIGHT_GRAPH[4004], RIGHT_GRAPH[3940], RIGHT_GRAPH[3876], RIGHT_GRAPH[3812], RIGHT_GRAPH[3748], RIGHT_GRAPH[3684], RIGHT_GRAPH[3620]};
					9'd485	:	PATTERN = {RIGHT_GRAPH[4069], RIGHT_GRAPH[4005], RIGHT_GRAPH[3941], RIGHT_GRAPH[3877], RIGHT_GRAPH[3813], RIGHT_GRAPH[3749], RIGHT_GRAPH[3685], RIGHT_GRAPH[3621]};
					9'd486	:	PATTERN = {RIGHT_GRAPH[4070], RIGHT_GRAPH[4006], RIGHT_GRAPH[3942], RIGHT_GRAPH[3878], RIGHT_GRAPH[3814], RIGHT_GRAPH[3750], RIGHT_GRAPH[3686], RIGHT_GRAPH[3622]};
					9'd487	:	PATTERN = {RIGHT_GRAPH[4071], RIGHT_GRAPH[4007], RIGHT_GRAPH[3943], RIGHT_GRAPH[3879], RIGHT_GRAPH[3815], RIGHT_GRAPH[3751], RIGHT_GRAPH[3687], RIGHT_GRAPH[3623]};
					9'd488	:	PATTERN = {RIGHT_GRAPH[4072], RIGHT_GRAPH[4008], RIGHT_GRAPH[3944], RIGHT_GRAPH[3880], RIGHT_GRAPH[3816], RIGHT_GRAPH[3752], RIGHT_GRAPH[3688], RIGHT_GRAPH[3624]};
					9'd489	:	PATTERN = {RIGHT_GRAPH[4073], RIGHT_GRAPH[4009], RIGHT_GRAPH[3945], RIGHT_GRAPH[3881], RIGHT_GRAPH[3817], RIGHT_GRAPH[3753], RIGHT_GRAPH[3689], RIGHT_GRAPH[3625]};
					9'd490	:	PATTERN = {RIGHT_GRAPH[4074], RIGHT_GRAPH[4010], RIGHT_GRAPH[3946], RIGHT_GRAPH[3882], RIGHT_GRAPH[3818], RIGHT_GRAPH[3754], RIGHT_GRAPH[3690], RIGHT_GRAPH[3626]};
					9'd491	:	PATTERN = {RIGHT_GRAPH[4075], RIGHT_GRAPH[4011], RIGHT_GRAPH[3947], RIGHT_GRAPH[3883], RIGHT_GRAPH[3819], RIGHT_GRAPH[3755], RIGHT_GRAPH[3691], RIGHT_GRAPH[3627]};
					9'd492	:	PATTERN = {RIGHT_GRAPH[4076], RIGHT_GRAPH[4012], RIGHT_GRAPH[3948], RIGHT_GRAPH[3884], RIGHT_GRAPH[3820], RIGHT_GRAPH[3756], RIGHT_GRAPH[3692], RIGHT_GRAPH[3628]};
					9'd493	:	PATTERN = {RIGHT_GRAPH[4077], RIGHT_GRAPH[4013], RIGHT_GRAPH[3949], RIGHT_GRAPH[3885], RIGHT_GRAPH[3821], RIGHT_GRAPH[3757], RIGHT_GRAPH[3693], RIGHT_GRAPH[3629]};
					9'd494	:	PATTERN = {RIGHT_GRAPH[4078], RIGHT_GRAPH[4014], RIGHT_GRAPH[3950], RIGHT_GRAPH[3886], RIGHT_GRAPH[3822], RIGHT_GRAPH[3758], RIGHT_GRAPH[3694], RIGHT_GRAPH[3630]};
					9'd495	:	PATTERN = {RIGHT_GRAPH[4079], RIGHT_GRAPH[4015], RIGHT_GRAPH[3951], RIGHT_GRAPH[3887], RIGHT_GRAPH[3823], RIGHT_GRAPH[3759], RIGHT_GRAPH[3695], RIGHT_GRAPH[3631]};
					9'd496	:	PATTERN = {RIGHT_GRAPH[4080], RIGHT_GRAPH[4016], RIGHT_GRAPH[3952], RIGHT_GRAPH[3888], RIGHT_GRAPH[3824], RIGHT_GRAPH[3760], RIGHT_GRAPH[3696], RIGHT_GRAPH[3632]};
					9'd497	:	PATTERN = {RIGHT_GRAPH[4081], RIGHT_GRAPH[4017], RIGHT_GRAPH[3953], RIGHT_GRAPH[3889], RIGHT_GRAPH[3825], RIGHT_GRAPH[3761], RIGHT_GRAPH[3697], RIGHT_GRAPH[3633]};
					9'd498	:	PATTERN = {RIGHT_GRAPH[4082], RIGHT_GRAPH[4018], RIGHT_GRAPH[3954], RIGHT_GRAPH[3890], RIGHT_GRAPH[3826], RIGHT_GRAPH[3762], RIGHT_GRAPH[3698], RIGHT_GRAPH[3634]};
					9'd499	:	PATTERN = {RIGHT_GRAPH[4083], RIGHT_GRAPH[4019], RIGHT_GRAPH[3955], RIGHT_GRAPH[3891], RIGHT_GRAPH[3827], RIGHT_GRAPH[3763], RIGHT_GRAPH[3699], RIGHT_GRAPH[3635]};
					9'd500	:	PATTERN = {RIGHT_GRAPH[4084], RIGHT_GRAPH[4020], RIGHT_GRAPH[3956], RIGHT_GRAPH[3892], RIGHT_GRAPH[3828], RIGHT_GRAPH[3764], RIGHT_GRAPH[3700], RIGHT_GRAPH[3636]};
					9'd501	:	PATTERN = {RIGHT_GRAPH[4085], RIGHT_GRAPH[4021], RIGHT_GRAPH[3957], RIGHT_GRAPH[3893], RIGHT_GRAPH[3829], RIGHT_GRAPH[3765], RIGHT_GRAPH[3701], RIGHT_GRAPH[3637]};
					9'd502	:	PATTERN = {RIGHT_GRAPH[4086], RIGHT_GRAPH[4022], RIGHT_GRAPH[3958], RIGHT_GRAPH[3894], RIGHT_GRAPH[3830], RIGHT_GRAPH[3766], RIGHT_GRAPH[3702], RIGHT_GRAPH[3638]};
					9'd503	:	PATTERN = {RIGHT_GRAPH[4087], RIGHT_GRAPH[4023], RIGHT_GRAPH[3959], RIGHT_GRAPH[3895], RIGHT_GRAPH[3831], RIGHT_GRAPH[3767], RIGHT_GRAPH[3703], RIGHT_GRAPH[3639]};
					9'd504	:	PATTERN = {RIGHT_GRAPH[4088], RIGHT_GRAPH[4024], RIGHT_GRAPH[3960], RIGHT_GRAPH[3896], RIGHT_GRAPH[3832], RIGHT_GRAPH[3768], RIGHT_GRAPH[3704], RIGHT_GRAPH[3640]};
					9'd505	:	PATTERN = {RIGHT_GRAPH[4089], RIGHT_GRAPH[4025], RIGHT_GRAPH[3961], RIGHT_GRAPH[3897], RIGHT_GRAPH[3833], RIGHT_GRAPH[3769], RIGHT_GRAPH[3705], RIGHT_GRAPH[3641]};
					9'd506	:	PATTERN = {RIGHT_GRAPH[4090], RIGHT_GRAPH[4026], RIGHT_GRAPH[3962], RIGHT_GRAPH[3898], RIGHT_GRAPH[3834], RIGHT_GRAPH[3770], RIGHT_GRAPH[3706], RIGHT_GRAPH[3642]};
					9'd507	:	PATTERN = {RIGHT_GRAPH[4091], RIGHT_GRAPH[4027], RIGHT_GRAPH[3963], RIGHT_GRAPH[3899], RIGHT_GRAPH[3835], RIGHT_GRAPH[3771], RIGHT_GRAPH[3707], RIGHT_GRAPH[3643]};
					9'd508	:	PATTERN = {RIGHT_GRAPH[4092], RIGHT_GRAPH[4028], RIGHT_GRAPH[3964], RIGHT_GRAPH[3900], RIGHT_GRAPH[3836], RIGHT_GRAPH[3772], RIGHT_GRAPH[3708], RIGHT_GRAPH[3644]};
					9'd509	:	PATTERN = {RIGHT_GRAPH[4093], RIGHT_GRAPH[4029], RIGHT_GRAPH[3965], RIGHT_GRAPH[3901], RIGHT_GRAPH[3837], RIGHT_GRAPH[3773], RIGHT_GRAPH[3709], RIGHT_GRAPH[3645]};
					9'd510	:	PATTERN = {RIGHT_GRAPH[4094], RIGHT_GRAPH[4030], RIGHT_GRAPH[3966], RIGHT_GRAPH[3902], RIGHT_GRAPH[3838], RIGHT_GRAPH[3774], RIGHT_GRAPH[3710], RIGHT_GRAPH[3646]};
					9'd511	:	PATTERN = {RIGHT_GRAPH[4095], RIGHT_GRAPH[4031], RIGHT_GRAPH[3967], RIGHT_GRAPH[3903], RIGHT_GRAPH[3839], RIGHT_GRAPH[3775], RIGHT_GRAPH[3711], RIGHT_GRAPH[3647]};		  
				endcase
			1'b1:
				case (INDEX)
				//------PAGE 0-------//
				  	9'd  0	:	PATTERN = {LEFT_GRAPH[ 448], LEFT_GRAPH[ 384], LEFT_GRAPH[ 320], LEFT_GRAPH[ 256], LEFT_GRAPH[ 192], LEFT_GRAPH[ 128], LEFT_GRAPH[  64], LEFT_GRAPH[   0]};
					9'd  1	:	PATTERN = {LEFT_GRAPH[ 449], LEFT_GRAPH[ 385], LEFT_GRAPH[ 321], LEFT_GRAPH[ 257], LEFT_GRAPH[ 193], LEFT_GRAPH[ 129], LEFT_GRAPH[  65], LEFT_GRAPH[   1]};
					9'd  2	:	PATTERN = {LEFT_GRAPH[ 450], LEFT_GRAPH[ 386], LEFT_GRAPH[ 322], LEFT_GRAPH[ 258], LEFT_GRAPH[ 194], LEFT_GRAPH[ 130], LEFT_GRAPH[  66], LEFT_GRAPH[   2]};
					9'd  3	:	PATTERN = {LEFT_GRAPH[ 451], LEFT_GRAPH[ 387], LEFT_GRAPH[ 323], LEFT_GRAPH[ 259], LEFT_GRAPH[ 195], LEFT_GRAPH[ 131], LEFT_GRAPH[  67], LEFT_GRAPH[   3]};
					9'd  4	:	PATTERN = {LEFT_GRAPH[ 452], LEFT_GRAPH[ 388], LEFT_GRAPH[ 324], LEFT_GRAPH[ 260], LEFT_GRAPH[ 196], LEFT_GRAPH[ 132], LEFT_GRAPH[  68], LEFT_GRAPH[   4]};
					9'd  5	:	PATTERN = {LEFT_GRAPH[ 453], LEFT_GRAPH[ 389], LEFT_GRAPH[ 325], LEFT_GRAPH[ 261], LEFT_GRAPH[ 197], LEFT_GRAPH[ 133], LEFT_GRAPH[  69], LEFT_GRAPH[   5]};
					9'd  6	:	PATTERN = {LEFT_GRAPH[ 454], LEFT_GRAPH[ 390], LEFT_GRAPH[ 326], LEFT_GRAPH[ 262], LEFT_GRAPH[ 198], LEFT_GRAPH[ 134], LEFT_GRAPH[  70], LEFT_GRAPH[   6]};
					9'd  7	:	PATTERN = {LEFT_GRAPH[ 455], LEFT_GRAPH[ 391], LEFT_GRAPH[ 327], LEFT_GRAPH[ 263], LEFT_GRAPH[ 199], LEFT_GRAPH[ 135], LEFT_GRAPH[  71], LEFT_GRAPH[   7]};
					9'd  8	:	PATTERN = {LEFT_GRAPH[ 456], LEFT_GRAPH[ 392], LEFT_GRAPH[ 328], LEFT_GRAPH[ 264], LEFT_GRAPH[ 200], LEFT_GRAPH[ 136], LEFT_GRAPH[  72], LEFT_GRAPH[   8]};
					9'd  9	:	PATTERN = {LEFT_GRAPH[ 457], LEFT_GRAPH[ 393], LEFT_GRAPH[ 329], LEFT_GRAPH[ 265], LEFT_GRAPH[ 201], LEFT_GRAPH[ 137], LEFT_GRAPH[  73], LEFT_GRAPH[   9]};
					9'd 10	:	PATTERN = {LEFT_GRAPH[ 458], LEFT_GRAPH[ 394], LEFT_GRAPH[ 330], LEFT_GRAPH[ 266], LEFT_GRAPH[ 202], LEFT_GRAPH[ 138], LEFT_GRAPH[  74], LEFT_GRAPH[  10]};
					9'd 11	:	PATTERN = {LEFT_GRAPH[ 459], LEFT_GRAPH[ 395], LEFT_GRAPH[ 331], LEFT_GRAPH[ 267], LEFT_GRAPH[ 203], LEFT_GRAPH[ 139], LEFT_GRAPH[  75], LEFT_GRAPH[  11]};
					9'd 12	:	PATTERN = {LEFT_GRAPH[ 460], LEFT_GRAPH[ 396], LEFT_GRAPH[ 332], LEFT_GRAPH[ 268], LEFT_GRAPH[ 204], LEFT_GRAPH[ 140], LEFT_GRAPH[  76], LEFT_GRAPH[  12]};
					9'd 13	:	PATTERN = {LEFT_GRAPH[ 461], LEFT_GRAPH[ 397], LEFT_GRAPH[ 333], LEFT_GRAPH[ 269], LEFT_GRAPH[ 205], LEFT_GRAPH[ 141], LEFT_GRAPH[  77], LEFT_GRAPH[  13]};
					9'd 14	:	PATTERN = {LEFT_GRAPH[ 462], LEFT_GRAPH[ 398], LEFT_GRAPH[ 334], LEFT_GRAPH[ 270], LEFT_GRAPH[ 206], LEFT_GRAPH[ 142], LEFT_GRAPH[  78], LEFT_GRAPH[  14]};
					9'd 15	:	PATTERN = {LEFT_GRAPH[ 463], LEFT_GRAPH[ 399], LEFT_GRAPH[ 335], LEFT_GRAPH[ 271], LEFT_GRAPH[ 207], LEFT_GRAPH[ 143], LEFT_GRAPH[  79], LEFT_GRAPH[  15]};
					9'd 16	:	PATTERN = {LEFT_GRAPH[ 464], LEFT_GRAPH[ 400], LEFT_GRAPH[ 336], LEFT_GRAPH[ 272], LEFT_GRAPH[ 208], LEFT_GRAPH[ 144], LEFT_GRAPH[  80], LEFT_GRAPH[  16]};
					9'd 17	:	PATTERN = {LEFT_GRAPH[ 465], LEFT_GRAPH[ 401], LEFT_GRAPH[ 337], LEFT_GRAPH[ 273], LEFT_GRAPH[ 209], LEFT_GRAPH[ 145], LEFT_GRAPH[  81], LEFT_GRAPH[  17]};
					9'd 18	:	PATTERN = {LEFT_GRAPH[ 466], LEFT_GRAPH[ 402], LEFT_GRAPH[ 338], LEFT_GRAPH[ 274], LEFT_GRAPH[ 210], LEFT_GRAPH[ 146], LEFT_GRAPH[  82], LEFT_GRAPH[  18]};
					9'd 19	:	PATTERN = {LEFT_GRAPH[ 467], LEFT_GRAPH[ 403], LEFT_GRAPH[ 339], LEFT_GRAPH[ 275], LEFT_GRAPH[ 211], LEFT_GRAPH[ 147], LEFT_GRAPH[  83], LEFT_GRAPH[  19]};
					9'd 20	:	PATTERN = {LEFT_GRAPH[ 468], LEFT_GRAPH[ 404], LEFT_GRAPH[ 340], LEFT_GRAPH[ 276], LEFT_GRAPH[ 212], LEFT_GRAPH[ 148], LEFT_GRAPH[  84], LEFT_GRAPH[  20]};
					9'd 21	:	PATTERN = {LEFT_GRAPH[ 469], LEFT_GRAPH[ 405], LEFT_GRAPH[ 341], LEFT_GRAPH[ 277], LEFT_GRAPH[ 213], LEFT_GRAPH[ 149], LEFT_GRAPH[  85], LEFT_GRAPH[  21]};
					9'd 22	:	PATTERN = {LEFT_GRAPH[ 470], LEFT_GRAPH[ 406], LEFT_GRAPH[ 342], LEFT_GRAPH[ 278], LEFT_GRAPH[ 214], LEFT_GRAPH[ 150], LEFT_GRAPH[  86], LEFT_GRAPH[  22]};
					9'd 23	:	PATTERN = {LEFT_GRAPH[ 471], LEFT_GRAPH[ 407], LEFT_GRAPH[ 343], LEFT_GRAPH[ 279], LEFT_GRAPH[ 215], LEFT_GRAPH[ 151], LEFT_GRAPH[  87], LEFT_GRAPH[  23]};
					9'd 24	:	PATTERN = {LEFT_GRAPH[ 472], LEFT_GRAPH[ 408], LEFT_GRAPH[ 344], LEFT_GRAPH[ 280], LEFT_GRAPH[ 216], LEFT_GRAPH[ 152], LEFT_GRAPH[  88], LEFT_GRAPH[  24]};
					9'd 25	:	PATTERN = {LEFT_GRAPH[ 473], LEFT_GRAPH[ 409], LEFT_GRAPH[ 345], LEFT_GRAPH[ 281], LEFT_GRAPH[ 217], LEFT_GRAPH[ 153], LEFT_GRAPH[  89], LEFT_GRAPH[  25]};
					9'd 26	:	PATTERN = {LEFT_GRAPH[ 474], LEFT_GRAPH[ 410], LEFT_GRAPH[ 346], LEFT_GRAPH[ 282], LEFT_GRAPH[ 218], LEFT_GRAPH[ 154], LEFT_GRAPH[  90], LEFT_GRAPH[  26]};
					9'd 27	:	PATTERN = {LEFT_GRAPH[ 475], LEFT_GRAPH[ 411], LEFT_GRAPH[ 347], LEFT_GRAPH[ 283], LEFT_GRAPH[ 219], LEFT_GRAPH[ 155], LEFT_GRAPH[  91], LEFT_GRAPH[  27]};
					9'd 28	:	PATTERN = {LEFT_GRAPH[ 476], LEFT_GRAPH[ 412], LEFT_GRAPH[ 348], LEFT_GRAPH[ 284], LEFT_GRAPH[ 220], LEFT_GRAPH[ 156], LEFT_GRAPH[  92], LEFT_GRAPH[  28]};
					9'd 29	:	PATTERN = {LEFT_GRAPH[ 477], LEFT_GRAPH[ 413], LEFT_GRAPH[ 349], LEFT_GRAPH[ 285], LEFT_GRAPH[ 221], LEFT_GRAPH[ 157], LEFT_GRAPH[  93], LEFT_GRAPH[  29]};
					9'd 30	:	PATTERN = {LEFT_GRAPH[ 478], LEFT_GRAPH[ 414], LEFT_GRAPH[ 350], LEFT_GRAPH[ 286], LEFT_GRAPH[ 222], LEFT_GRAPH[ 158], LEFT_GRAPH[  94], LEFT_GRAPH[  30]};
					9'd 31	:	PATTERN = {LEFT_GRAPH[ 479], LEFT_GRAPH[ 415], LEFT_GRAPH[ 351], LEFT_GRAPH[ 287], LEFT_GRAPH[ 223], LEFT_GRAPH[ 159], LEFT_GRAPH[  95], LEFT_GRAPH[  31]};
					9'd 32	:	PATTERN = {LEFT_GRAPH[ 480], LEFT_GRAPH[ 416], LEFT_GRAPH[ 352], LEFT_GRAPH[ 288], LEFT_GRAPH[ 224], LEFT_GRAPH[ 160], LEFT_GRAPH[  96], LEFT_GRAPH[  32]};
					9'd 33	:	PATTERN = {LEFT_GRAPH[ 481], LEFT_GRAPH[ 417], LEFT_GRAPH[ 353], LEFT_GRAPH[ 289], LEFT_GRAPH[ 225], LEFT_GRAPH[ 161], LEFT_GRAPH[  97], LEFT_GRAPH[  33]};
					9'd 34	:	PATTERN = {LEFT_GRAPH[ 482], LEFT_GRAPH[ 418], LEFT_GRAPH[ 354], LEFT_GRAPH[ 290], LEFT_GRAPH[ 226], LEFT_GRAPH[ 162], LEFT_GRAPH[  98], LEFT_GRAPH[  34]};
					9'd 35	:	PATTERN = {LEFT_GRAPH[ 483], LEFT_GRAPH[ 419], LEFT_GRAPH[ 355], LEFT_GRAPH[ 291], LEFT_GRAPH[ 227], LEFT_GRAPH[ 163], LEFT_GRAPH[  99], LEFT_GRAPH[  35]};
					9'd 36	:	PATTERN = {LEFT_GRAPH[ 484], LEFT_GRAPH[ 420], LEFT_GRAPH[ 356], LEFT_GRAPH[ 292], LEFT_GRAPH[ 228], LEFT_GRAPH[ 164], LEFT_GRAPH[ 100], LEFT_GRAPH[  36]};
					9'd 37	:	PATTERN = {LEFT_GRAPH[ 485], LEFT_GRAPH[ 421], LEFT_GRAPH[ 357], LEFT_GRAPH[ 293], LEFT_GRAPH[ 229], LEFT_GRAPH[ 165], LEFT_GRAPH[ 101], LEFT_GRAPH[  37]};
					9'd 38	:	PATTERN = {LEFT_GRAPH[ 486], LEFT_GRAPH[ 422], LEFT_GRAPH[ 358], LEFT_GRAPH[ 294], LEFT_GRAPH[ 230], LEFT_GRAPH[ 166], LEFT_GRAPH[ 102], LEFT_GRAPH[  38]};
					9'd 39	:	PATTERN = {LEFT_GRAPH[ 487], LEFT_GRAPH[ 423], LEFT_GRAPH[ 359], LEFT_GRAPH[ 295], LEFT_GRAPH[ 231], LEFT_GRAPH[ 167], LEFT_GRAPH[ 103], LEFT_GRAPH[  39]};
					9'd 40	:	PATTERN = {LEFT_GRAPH[ 488], LEFT_GRAPH[ 424], LEFT_GRAPH[ 360], LEFT_GRAPH[ 296], LEFT_GRAPH[ 232], LEFT_GRAPH[ 168], LEFT_GRAPH[ 104], LEFT_GRAPH[  40]};
					9'd 41	:	PATTERN = {LEFT_GRAPH[ 489], LEFT_GRAPH[ 425], LEFT_GRAPH[ 361], LEFT_GRAPH[ 297], LEFT_GRAPH[ 233], LEFT_GRAPH[ 169], LEFT_GRAPH[ 105], LEFT_GRAPH[  41]};
					9'd 42	:	PATTERN = {LEFT_GRAPH[ 490], LEFT_GRAPH[ 426], LEFT_GRAPH[ 362], LEFT_GRAPH[ 298], LEFT_GRAPH[ 234], LEFT_GRAPH[ 170], LEFT_GRAPH[ 106], LEFT_GRAPH[  42]};
					9'd 43	:	PATTERN = {LEFT_GRAPH[ 491], LEFT_GRAPH[ 427], LEFT_GRAPH[ 363], LEFT_GRAPH[ 299], LEFT_GRAPH[ 235], LEFT_GRAPH[ 171], LEFT_GRAPH[ 107], LEFT_GRAPH[  43]};
					9'd 44	:	PATTERN = {LEFT_GRAPH[ 492], LEFT_GRAPH[ 428], LEFT_GRAPH[ 364], LEFT_GRAPH[ 300], LEFT_GRAPH[ 236], LEFT_GRAPH[ 172], LEFT_GRAPH[ 108], LEFT_GRAPH[  44]};
					9'd 45	:	PATTERN = {LEFT_GRAPH[ 493], LEFT_GRAPH[ 429], LEFT_GRAPH[ 365], LEFT_GRAPH[ 301], LEFT_GRAPH[ 237], LEFT_GRAPH[ 173], LEFT_GRAPH[ 109], LEFT_GRAPH[  45]};
					9'd 46	:	PATTERN = {LEFT_GRAPH[ 494], LEFT_GRAPH[ 430], LEFT_GRAPH[ 366], LEFT_GRAPH[ 302], LEFT_GRAPH[ 238], LEFT_GRAPH[ 174], LEFT_GRAPH[ 110], LEFT_GRAPH[  46]};
					9'd 47	:	PATTERN = {LEFT_GRAPH[ 495], LEFT_GRAPH[ 431], LEFT_GRAPH[ 367], LEFT_GRAPH[ 303], LEFT_GRAPH[ 239], LEFT_GRAPH[ 175], LEFT_GRAPH[ 111], LEFT_GRAPH[  47]};
					9'd 48	:	PATTERN = {LEFT_GRAPH[ 496], LEFT_GRAPH[ 432], LEFT_GRAPH[ 368], LEFT_GRAPH[ 304], LEFT_GRAPH[ 240], LEFT_GRAPH[ 176], LEFT_GRAPH[ 112], LEFT_GRAPH[  48]};
					9'd 49	:	PATTERN = {LEFT_GRAPH[ 497], LEFT_GRAPH[ 433], LEFT_GRAPH[ 369], LEFT_GRAPH[ 305], LEFT_GRAPH[ 241], LEFT_GRAPH[ 177], LEFT_GRAPH[ 113], LEFT_GRAPH[  49]};
					9'd 50	:	PATTERN = {LEFT_GRAPH[ 498], LEFT_GRAPH[ 434], LEFT_GRAPH[ 370], LEFT_GRAPH[ 306], LEFT_GRAPH[ 242], LEFT_GRAPH[ 178], LEFT_GRAPH[ 114], LEFT_GRAPH[  50]};
					9'd 51	:	PATTERN = {LEFT_GRAPH[ 499], LEFT_GRAPH[ 435], LEFT_GRAPH[ 371], LEFT_GRAPH[ 307], LEFT_GRAPH[ 243], LEFT_GRAPH[ 179], LEFT_GRAPH[ 115], LEFT_GRAPH[  51]};
					9'd 52	:	PATTERN = {LEFT_GRAPH[ 500], LEFT_GRAPH[ 436], LEFT_GRAPH[ 372], LEFT_GRAPH[ 308], LEFT_GRAPH[ 244], LEFT_GRAPH[ 180], LEFT_GRAPH[ 116], LEFT_GRAPH[  52]};
					9'd 53	:	PATTERN = {LEFT_GRAPH[ 501], LEFT_GRAPH[ 437], LEFT_GRAPH[ 373], LEFT_GRAPH[ 309], LEFT_GRAPH[ 245], LEFT_GRAPH[ 181], LEFT_GRAPH[ 117], LEFT_GRAPH[  53]};
					9'd 54	:	PATTERN = {LEFT_GRAPH[ 502], LEFT_GRAPH[ 438], LEFT_GRAPH[ 374], LEFT_GRAPH[ 310], LEFT_GRAPH[ 246], LEFT_GRAPH[ 182], LEFT_GRAPH[ 118], LEFT_GRAPH[  54]};
					9'd 55	:	PATTERN = {LEFT_GRAPH[ 503], LEFT_GRAPH[ 439], LEFT_GRAPH[ 375], LEFT_GRAPH[ 311], LEFT_GRAPH[ 247], LEFT_GRAPH[ 183], LEFT_GRAPH[ 119], LEFT_GRAPH[  55]};
					9'd 56	:	PATTERN = {LEFT_GRAPH[ 504], LEFT_GRAPH[ 440], LEFT_GRAPH[ 376], LEFT_GRAPH[ 312], LEFT_GRAPH[ 248], LEFT_GRAPH[ 184], LEFT_GRAPH[ 120], LEFT_GRAPH[  56]};
					9'd 57	:	PATTERN = {LEFT_GRAPH[ 505], LEFT_GRAPH[ 441], LEFT_GRAPH[ 377], LEFT_GRAPH[ 313], LEFT_GRAPH[ 249], LEFT_GRAPH[ 185], LEFT_GRAPH[ 121], LEFT_GRAPH[  57]};
					9'd 58	:	PATTERN = {LEFT_GRAPH[ 506], LEFT_GRAPH[ 442], LEFT_GRAPH[ 378], LEFT_GRAPH[ 314], LEFT_GRAPH[ 250], LEFT_GRAPH[ 186], LEFT_GRAPH[ 122], LEFT_GRAPH[  58]};
					9'd 59	:	PATTERN = {LEFT_GRAPH[ 507], LEFT_GRAPH[ 443], LEFT_GRAPH[ 379], LEFT_GRAPH[ 315], LEFT_GRAPH[ 251], LEFT_GRAPH[ 187], LEFT_GRAPH[ 123], LEFT_GRAPH[  59]};
					9'd 60	:	PATTERN = {LEFT_GRAPH[ 508], LEFT_GRAPH[ 444], LEFT_GRAPH[ 380], LEFT_GRAPH[ 316], LEFT_GRAPH[ 252], LEFT_GRAPH[ 188], LEFT_GRAPH[ 124], LEFT_GRAPH[  60]};
					9'd 61	:	PATTERN = {LEFT_GRAPH[ 509], LEFT_GRAPH[ 445], LEFT_GRAPH[ 381], LEFT_GRAPH[ 317], LEFT_GRAPH[ 253], LEFT_GRAPH[ 189], LEFT_GRAPH[ 125], LEFT_GRAPH[  61]};
					9'd 62	:	PATTERN = {LEFT_GRAPH[ 510], LEFT_GRAPH[ 446], LEFT_GRAPH[ 382], LEFT_GRAPH[ 318], LEFT_GRAPH[ 254], LEFT_GRAPH[ 190], LEFT_GRAPH[ 126], LEFT_GRAPH[  62]};
					9'd 63	:	PATTERN = {LEFT_GRAPH[ 511], LEFT_GRAPH[ 447], LEFT_GRAPH[ 383], LEFT_GRAPH[ 319], LEFT_GRAPH[ 255], LEFT_GRAPH[ 191], LEFT_GRAPH[ 127], LEFT_GRAPH[  63]};
					9'd 64	:	PATTERN = {LEFT_GRAPH[ 960], LEFT_GRAPH[ 896], LEFT_GRAPH[ 832], LEFT_GRAPH[ 768], LEFT_GRAPH[ 704], LEFT_GRAPH[ 640], LEFT_GRAPH[ 576], LEFT_GRAPH[ 512]};
					9'd 65	:	PATTERN = {LEFT_GRAPH[ 961], LEFT_GRAPH[ 897], LEFT_GRAPH[ 833], LEFT_GRAPH[ 769], LEFT_GRAPH[ 705], LEFT_GRAPH[ 641], LEFT_GRAPH[ 577], LEFT_GRAPH[ 513]};
					9'd 66	:	PATTERN = {LEFT_GRAPH[ 962], LEFT_GRAPH[ 898], LEFT_GRAPH[ 834], LEFT_GRAPH[ 770], LEFT_GRAPH[ 706], LEFT_GRAPH[ 642], LEFT_GRAPH[ 578], LEFT_GRAPH[ 514]};
					9'd 67	:	PATTERN = {LEFT_GRAPH[ 963], LEFT_GRAPH[ 899], LEFT_GRAPH[ 835], LEFT_GRAPH[ 771], LEFT_GRAPH[ 707], LEFT_GRAPH[ 643], LEFT_GRAPH[ 579], LEFT_GRAPH[ 515]};
					9'd 68	:	PATTERN = {LEFT_GRAPH[ 964], LEFT_GRAPH[ 900], LEFT_GRAPH[ 836], LEFT_GRAPH[ 772], LEFT_GRAPH[ 708], LEFT_GRAPH[ 644], LEFT_GRAPH[ 580], LEFT_GRAPH[ 516]};
					9'd 69	:	PATTERN = {LEFT_GRAPH[ 965], LEFT_GRAPH[ 901], LEFT_GRAPH[ 837], LEFT_GRAPH[ 773], LEFT_GRAPH[ 709], LEFT_GRAPH[ 645], LEFT_GRAPH[ 581], LEFT_GRAPH[ 517]};
					9'd 70	:	PATTERN = {LEFT_GRAPH[ 966], LEFT_GRAPH[ 902], LEFT_GRAPH[ 838], LEFT_GRAPH[ 774], LEFT_GRAPH[ 710], LEFT_GRAPH[ 646], LEFT_GRAPH[ 582], LEFT_GRAPH[ 518]};
					9'd 71	:	PATTERN = {LEFT_GRAPH[ 967], LEFT_GRAPH[ 903], LEFT_GRAPH[ 839], LEFT_GRAPH[ 775], LEFT_GRAPH[ 711], LEFT_GRAPH[ 647], LEFT_GRAPH[ 583], LEFT_GRAPH[ 519]};
					9'd 72	:	PATTERN = {LEFT_GRAPH[ 968], LEFT_GRAPH[ 904], LEFT_GRAPH[ 840], LEFT_GRAPH[ 776], LEFT_GRAPH[ 712], LEFT_GRAPH[ 648], LEFT_GRAPH[ 584], LEFT_GRAPH[ 520]};
					9'd 73	:	PATTERN = {LEFT_GRAPH[ 969], LEFT_GRAPH[ 905], LEFT_GRAPH[ 841], LEFT_GRAPH[ 777], LEFT_GRAPH[ 713], LEFT_GRAPH[ 649], LEFT_GRAPH[ 585], LEFT_GRAPH[ 521]};
					9'd 74	:	PATTERN = {LEFT_GRAPH[ 970], LEFT_GRAPH[ 906], LEFT_GRAPH[ 842], LEFT_GRAPH[ 778], LEFT_GRAPH[ 714], LEFT_GRAPH[ 650], LEFT_GRAPH[ 586], LEFT_GRAPH[ 522]};
					9'd 75	:	PATTERN = {LEFT_GRAPH[ 971], LEFT_GRAPH[ 907], LEFT_GRAPH[ 843], LEFT_GRAPH[ 779], LEFT_GRAPH[ 715], LEFT_GRAPH[ 651], LEFT_GRAPH[ 587], LEFT_GRAPH[ 523]};
					9'd 76	:	PATTERN = {LEFT_GRAPH[ 972], LEFT_GRAPH[ 908], LEFT_GRAPH[ 844], LEFT_GRAPH[ 780], LEFT_GRAPH[ 716], LEFT_GRAPH[ 652], LEFT_GRAPH[ 588], LEFT_GRAPH[ 524]};
					9'd 77	:	PATTERN = {LEFT_GRAPH[ 973], LEFT_GRAPH[ 909], LEFT_GRAPH[ 845], LEFT_GRAPH[ 781], LEFT_GRAPH[ 717], LEFT_GRAPH[ 653], LEFT_GRAPH[ 589], LEFT_GRAPH[ 525]};
					9'd 78	:	PATTERN = {LEFT_GRAPH[ 974], LEFT_GRAPH[ 910], LEFT_GRAPH[ 846], LEFT_GRAPH[ 782], LEFT_GRAPH[ 718], LEFT_GRAPH[ 654], LEFT_GRAPH[ 590], LEFT_GRAPH[ 526]};
					9'd 79	:	PATTERN = {LEFT_GRAPH[ 975], LEFT_GRAPH[ 911], LEFT_GRAPH[ 847], LEFT_GRAPH[ 783], LEFT_GRAPH[ 719], LEFT_GRAPH[ 655], LEFT_GRAPH[ 591], LEFT_GRAPH[ 527]};
					9'd 80	:	PATTERN = {LEFT_GRAPH[ 976], LEFT_GRAPH[ 912], LEFT_GRAPH[ 848], LEFT_GRAPH[ 784], LEFT_GRAPH[ 720], LEFT_GRAPH[ 656], LEFT_GRAPH[ 592], LEFT_GRAPH[ 528]};
					9'd 81	:	PATTERN = {LEFT_GRAPH[ 977], LEFT_GRAPH[ 913], LEFT_GRAPH[ 849], LEFT_GRAPH[ 785], LEFT_GRAPH[ 721], LEFT_GRAPH[ 657], LEFT_GRAPH[ 593], LEFT_GRAPH[ 529]};
					9'd 82	:	PATTERN = {LEFT_GRAPH[ 978], LEFT_GRAPH[ 914], LEFT_GRAPH[ 850], LEFT_GRAPH[ 786], LEFT_GRAPH[ 722], LEFT_GRAPH[ 658], LEFT_GRAPH[ 594], LEFT_GRAPH[ 530]};
					9'd 83	:	PATTERN = {LEFT_GRAPH[ 979], LEFT_GRAPH[ 915], LEFT_GRAPH[ 851], LEFT_GRAPH[ 787], LEFT_GRAPH[ 723], LEFT_GRAPH[ 659], LEFT_GRAPH[ 595], LEFT_GRAPH[ 531]};
					9'd 84	:	PATTERN = {LEFT_GRAPH[ 980], LEFT_GRAPH[ 916], LEFT_GRAPH[ 852], LEFT_GRAPH[ 788], LEFT_GRAPH[ 724], LEFT_GRAPH[ 660], LEFT_GRAPH[ 596], LEFT_GRAPH[ 532]};
					9'd 85	:	PATTERN = {LEFT_GRAPH[ 981], LEFT_GRAPH[ 917], LEFT_GRAPH[ 853], LEFT_GRAPH[ 789], LEFT_GRAPH[ 725], LEFT_GRAPH[ 661], LEFT_GRAPH[ 597], LEFT_GRAPH[ 533]};
					9'd 86	:	PATTERN = {LEFT_GRAPH[ 982], LEFT_GRAPH[ 918], LEFT_GRAPH[ 854], LEFT_GRAPH[ 790], LEFT_GRAPH[ 726], LEFT_GRAPH[ 662], LEFT_GRAPH[ 598], LEFT_GRAPH[ 534]};
					9'd 87	:	PATTERN = {LEFT_GRAPH[ 983], LEFT_GRAPH[ 919], LEFT_GRAPH[ 855], LEFT_GRAPH[ 791], LEFT_GRAPH[ 727], LEFT_GRAPH[ 663], LEFT_GRAPH[ 599], LEFT_GRAPH[ 535]};
					9'd 88	:	PATTERN = {LEFT_GRAPH[ 984], LEFT_GRAPH[ 920], LEFT_GRAPH[ 856], LEFT_GRAPH[ 792], LEFT_GRAPH[ 728], LEFT_GRAPH[ 664], LEFT_GRAPH[ 600], LEFT_GRAPH[ 536]};
					9'd 89	:	PATTERN = {LEFT_GRAPH[ 985], LEFT_GRAPH[ 921], LEFT_GRAPH[ 857], LEFT_GRAPH[ 793], LEFT_GRAPH[ 729], LEFT_GRAPH[ 665], LEFT_GRAPH[ 601], LEFT_GRAPH[ 537]};
					9'd 90	:	PATTERN = {LEFT_GRAPH[ 986], LEFT_GRAPH[ 922], LEFT_GRAPH[ 858], LEFT_GRAPH[ 794], LEFT_GRAPH[ 730], LEFT_GRAPH[ 666], LEFT_GRAPH[ 602], LEFT_GRAPH[ 538]};
					9'd 91	:	PATTERN = {LEFT_GRAPH[ 987], LEFT_GRAPH[ 923], LEFT_GRAPH[ 859], LEFT_GRAPH[ 795], LEFT_GRAPH[ 731], LEFT_GRAPH[ 667], LEFT_GRAPH[ 603], LEFT_GRAPH[ 539]};
					9'd 92	:	PATTERN = {LEFT_GRAPH[ 988], LEFT_GRAPH[ 924], LEFT_GRAPH[ 860], LEFT_GRAPH[ 796], LEFT_GRAPH[ 732], LEFT_GRAPH[ 668], LEFT_GRAPH[ 604], LEFT_GRAPH[ 540]};
					9'd 93	:	PATTERN = {LEFT_GRAPH[ 989], LEFT_GRAPH[ 925], LEFT_GRAPH[ 861], LEFT_GRAPH[ 797], LEFT_GRAPH[ 733], LEFT_GRAPH[ 669], LEFT_GRAPH[ 605], LEFT_GRAPH[ 541]};
					9'd 94	:	PATTERN = {LEFT_GRAPH[ 990], LEFT_GRAPH[ 926], LEFT_GRAPH[ 862], LEFT_GRAPH[ 798], LEFT_GRAPH[ 734], LEFT_GRAPH[ 670], LEFT_GRAPH[ 606], LEFT_GRAPH[ 542]};
					9'd 95	:	PATTERN = {LEFT_GRAPH[ 991], LEFT_GRAPH[ 927], LEFT_GRAPH[ 863], LEFT_GRAPH[ 799], LEFT_GRAPH[ 735], LEFT_GRAPH[ 671], LEFT_GRAPH[ 607], LEFT_GRAPH[ 543]};
					9'd 96	:	PATTERN = {LEFT_GRAPH[ 992], LEFT_GRAPH[ 928], LEFT_GRAPH[ 864], LEFT_GRAPH[ 800], LEFT_GRAPH[ 736], LEFT_GRAPH[ 672], LEFT_GRAPH[ 608], LEFT_GRAPH[ 544]};
					9'd 97	:	PATTERN = {LEFT_GRAPH[ 993], LEFT_GRAPH[ 929], LEFT_GRAPH[ 865], LEFT_GRAPH[ 801], LEFT_GRAPH[ 737], LEFT_GRAPH[ 673], LEFT_GRAPH[ 609], LEFT_GRAPH[ 545]};
					9'd 98	:	PATTERN = {LEFT_GRAPH[ 994], LEFT_GRAPH[ 930], LEFT_GRAPH[ 866], LEFT_GRAPH[ 802], LEFT_GRAPH[ 738], LEFT_GRAPH[ 674], LEFT_GRAPH[ 610], LEFT_GRAPH[ 546]};
					9'd 99	:	PATTERN = {LEFT_GRAPH[ 995], LEFT_GRAPH[ 931], LEFT_GRAPH[ 867], LEFT_GRAPH[ 803], LEFT_GRAPH[ 739], LEFT_GRAPH[ 675], LEFT_GRAPH[ 611], LEFT_GRAPH[ 547]};
					9'd100	:	PATTERN = {LEFT_GRAPH[ 996], LEFT_GRAPH[ 932], LEFT_GRAPH[ 868], LEFT_GRAPH[ 804], LEFT_GRAPH[ 740], LEFT_GRAPH[ 676], LEFT_GRAPH[ 612], LEFT_GRAPH[ 548]};
					9'd101	:	PATTERN = {LEFT_GRAPH[ 997], LEFT_GRAPH[ 933], LEFT_GRAPH[ 869], LEFT_GRAPH[ 805], LEFT_GRAPH[ 741], LEFT_GRAPH[ 677], LEFT_GRAPH[ 613], LEFT_GRAPH[ 549]};
					9'd102	:	PATTERN = {LEFT_GRAPH[ 998], LEFT_GRAPH[ 934], LEFT_GRAPH[ 870], LEFT_GRAPH[ 806], LEFT_GRAPH[ 742], LEFT_GRAPH[ 678], LEFT_GRAPH[ 614], LEFT_GRAPH[ 550]};
					9'd103	:	PATTERN = {LEFT_GRAPH[ 999], LEFT_GRAPH[ 935], LEFT_GRAPH[ 871], LEFT_GRAPH[ 807], LEFT_GRAPH[ 743], LEFT_GRAPH[ 679], LEFT_GRAPH[ 615], LEFT_GRAPH[ 551]};
					9'd104	:	PATTERN = {LEFT_GRAPH[1000], LEFT_GRAPH[ 936], LEFT_GRAPH[ 872], LEFT_GRAPH[ 808], LEFT_GRAPH[ 744], LEFT_GRAPH[ 680], LEFT_GRAPH[ 616], LEFT_GRAPH[ 552]};
					9'd105	:	PATTERN = {LEFT_GRAPH[1001], LEFT_GRAPH[ 937], LEFT_GRAPH[ 873], LEFT_GRAPH[ 809], LEFT_GRAPH[ 745], LEFT_GRAPH[ 681], LEFT_GRAPH[ 617], LEFT_GRAPH[ 553]};
					9'd106	:	PATTERN = {LEFT_GRAPH[1002], LEFT_GRAPH[ 938], LEFT_GRAPH[ 874], LEFT_GRAPH[ 810], LEFT_GRAPH[ 746], LEFT_GRAPH[ 682], LEFT_GRAPH[ 618], LEFT_GRAPH[ 554]};
					9'd107	:	PATTERN = {LEFT_GRAPH[1003], LEFT_GRAPH[ 939], LEFT_GRAPH[ 875], LEFT_GRAPH[ 811], LEFT_GRAPH[ 747], LEFT_GRAPH[ 683], LEFT_GRAPH[ 619], LEFT_GRAPH[ 555]};
					9'd108	:	PATTERN = {LEFT_GRAPH[1004], LEFT_GRAPH[ 940], LEFT_GRAPH[ 876], LEFT_GRAPH[ 812], LEFT_GRAPH[ 748], LEFT_GRAPH[ 684], LEFT_GRAPH[ 620], LEFT_GRAPH[ 556]};
					9'd109	:	PATTERN = {LEFT_GRAPH[1005], LEFT_GRAPH[ 941], LEFT_GRAPH[ 877], LEFT_GRAPH[ 813], LEFT_GRAPH[ 749], LEFT_GRAPH[ 685], LEFT_GRAPH[ 621], LEFT_GRAPH[ 557]};
					9'd110	:	PATTERN = {LEFT_GRAPH[1006], LEFT_GRAPH[ 942], LEFT_GRAPH[ 878], LEFT_GRAPH[ 814], LEFT_GRAPH[ 750], LEFT_GRAPH[ 686], LEFT_GRAPH[ 622], LEFT_GRAPH[ 558]};
					9'd111	:	PATTERN = {LEFT_GRAPH[1007], LEFT_GRAPH[ 943], LEFT_GRAPH[ 879], LEFT_GRAPH[ 815], LEFT_GRAPH[ 751], LEFT_GRAPH[ 687], LEFT_GRAPH[ 623], LEFT_GRAPH[ 559]};
					9'd112	:	PATTERN = {LEFT_GRAPH[1008], LEFT_GRAPH[ 944], LEFT_GRAPH[ 880], LEFT_GRAPH[ 816], LEFT_GRAPH[ 752], LEFT_GRAPH[ 688], LEFT_GRAPH[ 624], LEFT_GRAPH[ 560]};
					9'd113	:	PATTERN = {LEFT_GRAPH[1009], LEFT_GRAPH[ 945], LEFT_GRAPH[ 881], LEFT_GRAPH[ 817], LEFT_GRAPH[ 753], LEFT_GRAPH[ 689], LEFT_GRAPH[ 625], LEFT_GRAPH[ 561]};
					9'd114	:	PATTERN = {LEFT_GRAPH[1010], LEFT_GRAPH[ 946], LEFT_GRAPH[ 882], LEFT_GRAPH[ 818], LEFT_GRAPH[ 754], LEFT_GRAPH[ 690], LEFT_GRAPH[ 626], LEFT_GRAPH[ 562]};
					9'd115	:	PATTERN = {LEFT_GRAPH[1011], LEFT_GRAPH[ 947], LEFT_GRAPH[ 883], LEFT_GRAPH[ 819], LEFT_GRAPH[ 755], LEFT_GRAPH[ 691], LEFT_GRAPH[ 627], LEFT_GRAPH[ 563]};
					9'd116	:	PATTERN = {LEFT_GRAPH[1012], LEFT_GRAPH[ 948], LEFT_GRAPH[ 884], LEFT_GRAPH[ 820], LEFT_GRAPH[ 756], LEFT_GRAPH[ 692], LEFT_GRAPH[ 628], LEFT_GRAPH[ 564]};
					9'd117	:	PATTERN = {LEFT_GRAPH[1013], LEFT_GRAPH[ 949], LEFT_GRAPH[ 885], LEFT_GRAPH[ 821], LEFT_GRAPH[ 757], LEFT_GRAPH[ 693], LEFT_GRAPH[ 629], LEFT_GRAPH[ 565]};
					9'd118	:	PATTERN = {LEFT_GRAPH[1014], LEFT_GRAPH[ 950], LEFT_GRAPH[ 886], LEFT_GRAPH[ 822], LEFT_GRAPH[ 758], LEFT_GRAPH[ 694], LEFT_GRAPH[ 630], LEFT_GRAPH[ 566]};
					9'd119	:	PATTERN = {LEFT_GRAPH[1015], LEFT_GRAPH[ 951], LEFT_GRAPH[ 887], LEFT_GRAPH[ 823], LEFT_GRAPH[ 759], LEFT_GRAPH[ 695], LEFT_GRAPH[ 631], LEFT_GRAPH[ 567]};
					9'd120	:	PATTERN = {LEFT_GRAPH[1016], LEFT_GRAPH[ 952], LEFT_GRAPH[ 888], LEFT_GRAPH[ 824], LEFT_GRAPH[ 760], LEFT_GRAPH[ 696], LEFT_GRAPH[ 632], LEFT_GRAPH[ 568]};
					9'd121	:	PATTERN = {LEFT_GRAPH[1017], LEFT_GRAPH[ 953], LEFT_GRAPH[ 889], LEFT_GRAPH[ 825], LEFT_GRAPH[ 761], LEFT_GRAPH[ 697], LEFT_GRAPH[ 633], LEFT_GRAPH[ 569]};
					9'd122	:	PATTERN = {LEFT_GRAPH[1018], LEFT_GRAPH[ 954], LEFT_GRAPH[ 890], LEFT_GRAPH[ 826], LEFT_GRAPH[ 762], LEFT_GRAPH[ 698], LEFT_GRAPH[ 634], LEFT_GRAPH[ 570]};
					9'd123	:	PATTERN = {LEFT_GRAPH[1019], LEFT_GRAPH[ 955], LEFT_GRAPH[ 891], LEFT_GRAPH[ 827], LEFT_GRAPH[ 763], LEFT_GRAPH[ 699], LEFT_GRAPH[ 635], LEFT_GRAPH[ 571]};
					9'd124	:	PATTERN = {LEFT_GRAPH[1020], LEFT_GRAPH[ 956], LEFT_GRAPH[ 892], LEFT_GRAPH[ 828], LEFT_GRAPH[ 764], LEFT_GRAPH[ 700], LEFT_GRAPH[ 636], LEFT_GRAPH[ 572]};
					9'd125	:	PATTERN = {LEFT_GRAPH[1021], LEFT_GRAPH[ 957], LEFT_GRAPH[ 893], LEFT_GRAPH[ 829], LEFT_GRAPH[ 765], LEFT_GRAPH[ 701], LEFT_GRAPH[ 637], LEFT_GRAPH[ 573]};
					9'd126	:	PATTERN = {LEFT_GRAPH[1022], LEFT_GRAPH[ 958], LEFT_GRAPH[ 894], LEFT_GRAPH[ 830], LEFT_GRAPH[ 766], LEFT_GRAPH[ 702], LEFT_GRAPH[ 638], LEFT_GRAPH[ 574]};
					9'd127	:	PATTERN = {LEFT_GRAPH[1023], LEFT_GRAPH[ 959], LEFT_GRAPH[ 895], LEFT_GRAPH[ 831], LEFT_GRAPH[ 767], LEFT_GRAPH[ 703], LEFT_GRAPH[ 639], LEFT_GRAPH[ 575]};
					9'd128	:	PATTERN = {LEFT_GRAPH[1472], LEFT_GRAPH[1408], LEFT_GRAPH[1344], LEFT_GRAPH[1280], LEFT_GRAPH[1216], LEFT_GRAPH[1152], LEFT_GRAPH[1088], LEFT_GRAPH[1024]};
					9'd129	:	PATTERN = {LEFT_GRAPH[1473], LEFT_GRAPH[1409], LEFT_GRAPH[1345], LEFT_GRAPH[1281], LEFT_GRAPH[1217], LEFT_GRAPH[1153], LEFT_GRAPH[1089], LEFT_GRAPH[1025]};
					9'd130	:	PATTERN = {LEFT_GRAPH[1474], LEFT_GRAPH[1410], LEFT_GRAPH[1346], LEFT_GRAPH[1282], LEFT_GRAPH[1218], LEFT_GRAPH[1154], LEFT_GRAPH[1090], LEFT_GRAPH[1026]};
					9'd131	:	PATTERN = {LEFT_GRAPH[1475], LEFT_GRAPH[1411], LEFT_GRAPH[1347], LEFT_GRAPH[1283], LEFT_GRAPH[1219], LEFT_GRAPH[1155], LEFT_GRAPH[1091], LEFT_GRAPH[1027]};
					9'd132	:	PATTERN = {LEFT_GRAPH[1476], LEFT_GRAPH[1412], LEFT_GRAPH[1348], LEFT_GRAPH[1284], LEFT_GRAPH[1220], LEFT_GRAPH[1156], LEFT_GRAPH[1092], LEFT_GRAPH[1028]};
					9'd133	:	PATTERN = {LEFT_GRAPH[1477], LEFT_GRAPH[1413], LEFT_GRAPH[1349], LEFT_GRAPH[1285], LEFT_GRAPH[1221], LEFT_GRAPH[1157], LEFT_GRAPH[1093], LEFT_GRAPH[1029]};
					9'd134	:	PATTERN = {LEFT_GRAPH[1478], LEFT_GRAPH[1414], LEFT_GRAPH[1350], LEFT_GRAPH[1286], LEFT_GRAPH[1222], LEFT_GRAPH[1158], LEFT_GRAPH[1094], LEFT_GRAPH[1030]};
					9'd135	:	PATTERN = {LEFT_GRAPH[1479], LEFT_GRAPH[1415], LEFT_GRAPH[1351], LEFT_GRAPH[1287], LEFT_GRAPH[1223], LEFT_GRAPH[1159], LEFT_GRAPH[1095], LEFT_GRAPH[1031]};
					9'd136	:	PATTERN = {LEFT_GRAPH[1480], LEFT_GRAPH[1416], LEFT_GRAPH[1352], LEFT_GRAPH[1288], LEFT_GRAPH[1224], LEFT_GRAPH[1160], LEFT_GRAPH[1096], LEFT_GRAPH[1032]};
					9'd137	:	PATTERN = {LEFT_GRAPH[1481], LEFT_GRAPH[1417], LEFT_GRAPH[1353], LEFT_GRAPH[1289], LEFT_GRAPH[1225], LEFT_GRAPH[1161], LEFT_GRAPH[1097], LEFT_GRAPH[1033]};
					9'd138	:	PATTERN = {LEFT_GRAPH[1482], LEFT_GRAPH[1418], LEFT_GRAPH[1354], LEFT_GRAPH[1290], LEFT_GRAPH[1226], LEFT_GRAPH[1162], LEFT_GRAPH[1098], LEFT_GRAPH[1034]};
					9'd139	:	PATTERN = {LEFT_GRAPH[1483], LEFT_GRAPH[1419], LEFT_GRAPH[1355], LEFT_GRAPH[1291], LEFT_GRAPH[1227], LEFT_GRAPH[1163], LEFT_GRAPH[1099], LEFT_GRAPH[1035]};
					9'd140	:	PATTERN = {LEFT_GRAPH[1484], LEFT_GRAPH[1420], LEFT_GRAPH[1356], LEFT_GRAPH[1292], LEFT_GRAPH[1228], LEFT_GRAPH[1164], LEFT_GRAPH[1100], LEFT_GRAPH[1036]};
					9'd141	:	PATTERN = {LEFT_GRAPH[1485], LEFT_GRAPH[1421], LEFT_GRAPH[1357], LEFT_GRAPH[1293], LEFT_GRAPH[1229], LEFT_GRAPH[1165], LEFT_GRAPH[1101], LEFT_GRAPH[1037]};
					9'd142	:	PATTERN = {LEFT_GRAPH[1486], LEFT_GRAPH[1422], LEFT_GRAPH[1358], LEFT_GRAPH[1294], LEFT_GRAPH[1230], LEFT_GRAPH[1166], LEFT_GRAPH[1102], LEFT_GRAPH[1038]};
					9'd143	:	PATTERN = {LEFT_GRAPH[1487], LEFT_GRAPH[1423], LEFT_GRAPH[1359], LEFT_GRAPH[1295], LEFT_GRAPH[1231], LEFT_GRAPH[1167], LEFT_GRAPH[1103], LEFT_GRAPH[1039]};
					9'd144	:	PATTERN = {LEFT_GRAPH[1488], LEFT_GRAPH[1424], LEFT_GRAPH[1360], LEFT_GRAPH[1296], LEFT_GRAPH[1232], LEFT_GRAPH[1168], LEFT_GRAPH[1104], LEFT_GRAPH[1040]};
					9'd145	:	PATTERN = {LEFT_GRAPH[1489], LEFT_GRAPH[1425], LEFT_GRAPH[1361], LEFT_GRAPH[1297], LEFT_GRAPH[1233], LEFT_GRAPH[1169], LEFT_GRAPH[1105], LEFT_GRAPH[1041]};
					9'd146	:	PATTERN = {LEFT_GRAPH[1490], LEFT_GRAPH[1426], LEFT_GRAPH[1362], LEFT_GRAPH[1298], LEFT_GRAPH[1234], LEFT_GRAPH[1170], LEFT_GRAPH[1106], LEFT_GRAPH[1042]};
					9'd147	:	PATTERN = {LEFT_GRAPH[1491], LEFT_GRAPH[1427], LEFT_GRAPH[1363], LEFT_GRAPH[1299], LEFT_GRAPH[1235], LEFT_GRAPH[1171], LEFT_GRAPH[1107], LEFT_GRAPH[1043]};
					9'd148	:	PATTERN = {LEFT_GRAPH[1492], LEFT_GRAPH[1428], LEFT_GRAPH[1364], LEFT_GRAPH[1300], LEFT_GRAPH[1236], LEFT_GRAPH[1172], LEFT_GRAPH[1108], LEFT_GRAPH[1044]};
					9'd149	:	PATTERN = {LEFT_GRAPH[1493], LEFT_GRAPH[1429], LEFT_GRAPH[1365], LEFT_GRAPH[1301], LEFT_GRAPH[1237], LEFT_GRAPH[1173], LEFT_GRAPH[1109], LEFT_GRAPH[1045]};
					9'd150	:	PATTERN = {LEFT_GRAPH[1494], LEFT_GRAPH[1430], LEFT_GRAPH[1366], LEFT_GRAPH[1302], LEFT_GRAPH[1238], LEFT_GRAPH[1174], LEFT_GRAPH[1110], LEFT_GRAPH[1046]};
					9'd151	:	PATTERN = {LEFT_GRAPH[1495], LEFT_GRAPH[1431], LEFT_GRAPH[1367], LEFT_GRAPH[1303], LEFT_GRAPH[1239], LEFT_GRAPH[1175], LEFT_GRAPH[1111], LEFT_GRAPH[1047]};
					9'd152	:	PATTERN = {LEFT_GRAPH[1496], LEFT_GRAPH[1432], LEFT_GRAPH[1368], LEFT_GRAPH[1304], LEFT_GRAPH[1240], LEFT_GRAPH[1176], LEFT_GRAPH[1112], LEFT_GRAPH[1048]};
					9'd153	:	PATTERN = {LEFT_GRAPH[1497], LEFT_GRAPH[1433], LEFT_GRAPH[1369], LEFT_GRAPH[1305], LEFT_GRAPH[1241], LEFT_GRAPH[1177], LEFT_GRAPH[1113], LEFT_GRAPH[1049]};
					9'd154	:	PATTERN = {LEFT_GRAPH[1498], LEFT_GRAPH[1434], LEFT_GRAPH[1370], LEFT_GRAPH[1306], LEFT_GRAPH[1242], LEFT_GRAPH[1178], LEFT_GRAPH[1114], LEFT_GRAPH[1050]};
					9'd155	:	PATTERN = {LEFT_GRAPH[1499], LEFT_GRAPH[1435], LEFT_GRAPH[1371], LEFT_GRAPH[1307], LEFT_GRAPH[1243], LEFT_GRAPH[1179], LEFT_GRAPH[1115], LEFT_GRAPH[1051]};
					9'd156	:	PATTERN = {LEFT_GRAPH[1500], LEFT_GRAPH[1436], LEFT_GRAPH[1372], LEFT_GRAPH[1308], LEFT_GRAPH[1244], LEFT_GRAPH[1180], LEFT_GRAPH[1116], LEFT_GRAPH[1052]};
					9'd157	:	PATTERN = {LEFT_GRAPH[1501], LEFT_GRAPH[1437], LEFT_GRAPH[1373], LEFT_GRAPH[1309], LEFT_GRAPH[1245], LEFT_GRAPH[1181], LEFT_GRAPH[1117], LEFT_GRAPH[1053]};
					9'd158	:	PATTERN = {LEFT_GRAPH[1502], LEFT_GRAPH[1438], LEFT_GRAPH[1374], LEFT_GRAPH[1310], LEFT_GRAPH[1246], LEFT_GRAPH[1182], LEFT_GRAPH[1118], LEFT_GRAPH[1054]};
					9'd159	:	PATTERN = {LEFT_GRAPH[1503], LEFT_GRAPH[1439], LEFT_GRAPH[1375], LEFT_GRAPH[1311], LEFT_GRAPH[1247], LEFT_GRAPH[1183], LEFT_GRAPH[1119], LEFT_GRAPH[1055]};
					9'd160	:	PATTERN = {LEFT_GRAPH[1504], LEFT_GRAPH[1440], LEFT_GRAPH[1376], LEFT_GRAPH[1312], LEFT_GRAPH[1248], LEFT_GRAPH[1184], LEFT_GRAPH[1120], LEFT_GRAPH[1056]};
					9'd161	:	PATTERN = {LEFT_GRAPH[1505], LEFT_GRAPH[1441], LEFT_GRAPH[1377], LEFT_GRAPH[1313], LEFT_GRAPH[1249], LEFT_GRAPH[1185], LEFT_GRAPH[1121], LEFT_GRAPH[1057]};
					9'd162	:	PATTERN = {LEFT_GRAPH[1506], LEFT_GRAPH[1442], LEFT_GRAPH[1378], LEFT_GRAPH[1314], LEFT_GRAPH[1250], LEFT_GRAPH[1186], LEFT_GRAPH[1122], LEFT_GRAPH[1058]};
					9'd163	:	PATTERN = {LEFT_GRAPH[1507], LEFT_GRAPH[1443], LEFT_GRAPH[1379], LEFT_GRAPH[1315], LEFT_GRAPH[1251], LEFT_GRAPH[1187], LEFT_GRAPH[1123], LEFT_GRAPH[1059]};
					9'd164	:	PATTERN = {LEFT_GRAPH[1508], LEFT_GRAPH[1444], LEFT_GRAPH[1380], LEFT_GRAPH[1316], LEFT_GRAPH[1252], LEFT_GRAPH[1188], LEFT_GRAPH[1124], LEFT_GRAPH[1060]};
					9'd165	:	PATTERN = {LEFT_GRAPH[1509], LEFT_GRAPH[1445], LEFT_GRAPH[1381], LEFT_GRAPH[1317], LEFT_GRAPH[1253], LEFT_GRAPH[1189], LEFT_GRAPH[1125], LEFT_GRAPH[1061]};
					9'd166	:	PATTERN = {LEFT_GRAPH[1510], LEFT_GRAPH[1446], LEFT_GRAPH[1382], LEFT_GRAPH[1318], LEFT_GRAPH[1254], LEFT_GRAPH[1190], LEFT_GRAPH[1126], LEFT_GRAPH[1062]};
					9'd167	:	PATTERN = {LEFT_GRAPH[1511], LEFT_GRAPH[1447], LEFT_GRAPH[1383], LEFT_GRAPH[1319], LEFT_GRAPH[1255], LEFT_GRAPH[1191], LEFT_GRAPH[1127], LEFT_GRAPH[1063]};
					9'd168	:	PATTERN = {LEFT_GRAPH[1512], LEFT_GRAPH[1448], LEFT_GRAPH[1384], LEFT_GRAPH[1320], LEFT_GRAPH[1256], LEFT_GRAPH[1192], LEFT_GRAPH[1128], LEFT_GRAPH[1064]};
					9'd169	:	PATTERN = {LEFT_GRAPH[1513], LEFT_GRAPH[1449], LEFT_GRAPH[1385], LEFT_GRAPH[1321], LEFT_GRAPH[1257], LEFT_GRAPH[1193], LEFT_GRAPH[1129], LEFT_GRAPH[1065]};
					9'd170	:	PATTERN = {LEFT_GRAPH[1514], LEFT_GRAPH[1450], LEFT_GRAPH[1386], LEFT_GRAPH[1322], LEFT_GRAPH[1258], LEFT_GRAPH[1194], LEFT_GRAPH[1130], LEFT_GRAPH[1066]};
					9'd171	:	PATTERN = {LEFT_GRAPH[1515], LEFT_GRAPH[1451], LEFT_GRAPH[1387], LEFT_GRAPH[1323], LEFT_GRAPH[1259], LEFT_GRAPH[1195], LEFT_GRAPH[1131], LEFT_GRAPH[1067]};
					9'd172	:	PATTERN = {LEFT_GRAPH[1516], LEFT_GRAPH[1452], LEFT_GRAPH[1388], LEFT_GRAPH[1324], LEFT_GRAPH[1260], LEFT_GRAPH[1196], LEFT_GRAPH[1132], LEFT_GRAPH[1068]};
					9'd173	:	PATTERN = {LEFT_GRAPH[1517], LEFT_GRAPH[1453], LEFT_GRAPH[1389], LEFT_GRAPH[1325], LEFT_GRAPH[1261], LEFT_GRAPH[1197], LEFT_GRAPH[1133], LEFT_GRAPH[1069]};
					9'd174	:	PATTERN = {LEFT_GRAPH[1518], LEFT_GRAPH[1454], LEFT_GRAPH[1390], LEFT_GRAPH[1326], LEFT_GRAPH[1262], LEFT_GRAPH[1198], LEFT_GRAPH[1134], LEFT_GRAPH[1070]};
					9'd175	:	PATTERN = {LEFT_GRAPH[1519], LEFT_GRAPH[1455], LEFT_GRAPH[1391], LEFT_GRAPH[1327], LEFT_GRAPH[1263], LEFT_GRAPH[1199], LEFT_GRAPH[1135], LEFT_GRAPH[1071]};
					9'd176	:	PATTERN = {LEFT_GRAPH[1520], LEFT_GRAPH[1456], LEFT_GRAPH[1392], LEFT_GRAPH[1328], LEFT_GRAPH[1264], LEFT_GRAPH[1200], LEFT_GRAPH[1136], LEFT_GRAPH[1072]};
					9'd177	:	PATTERN = {LEFT_GRAPH[1521], LEFT_GRAPH[1457], LEFT_GRAPH[1393], LEFT_GRAPH[1329], LEFT_GRAPH[1265], LEFT_GRAPH[1201], LEFT_GRAPH[1137], LEFT_GRAPH[1073]};
					9'd178	:	PATTERN = {LEFT_GRAPH[1522], LEFT_GRAPH[1458], LEFT_GRAPH[1394], LEFT_GRAPH[1330], LEFT_GRAPH[1266], LEFT_GRAPH[1202], LEFT_GRAPH[1138], LEFT_GRAPH[1074]};
					9'd179	:	PATTERN = {LEFT_GRAPH[1523], LEFT_GRAPH[1459], LEFT_GRAPH[1395], LEFT_GRAPH[1331], LEFT_GRAPH[1267], LEFT_GRAPH[1203], LEFT_GRAPH[1139], LEFT_GRAPH[1075]};
					9'd180	:	PATTERN = {LEFT_GRAPH[1524], LEFT_GRAPH[1460], LEFT_GRAPH[1396], LEFT_GRAPH[1332], LEFT_GRAPH[1268], LEFT_GRAPH[1204], LEFT_GRAPH[1140], LEFT_GRAPH[1076]};
					9'd181	:	PATTERN = {LEFT_GRAPH[1525], LEFT_GRAPH[1461], LEFT_GRAPH[1397], LEFT_GRAPH[1333], LEFT_GRAPH[1269], LEFT_GRAPH[1205], LEFT_GRAPH[1141], LEFT_GRAPH[1077]};
					9'd182	:	PATTERN = {LEFT_GRAPH[1526], LEFT_GRAPH[1462], LEFT_GRAPH[1398], LEFT_GRAPH[1334], LEFT_GRAPH[1270], LEFT_GRAPH[1206], LEFT_GRAPH[1142], LEFT_GRAPH[1078]};
					9'd183	:	PATTERN = {LEFT_GRAPH[1527], LEFT_GRAPH[1463], LEFT_GRAPH[1399], LEFT_GRAPH[1335], LEFT_GRAPH[1271], LEFT_GRAPH[1207], LEFT_GRAPH[1143], LEFT_GRAPH[1079]};
					9'd184	:	PATTERN = {LEFT_GRAPH[1528], LEFT_GRAPH[1464], LEFT_GRAPH[1400], LEFT_GRAPH[1336], LEFT_GRAPH[1272], LEFT_GRAPH[1208], LEFT_GRAPH[1144], LEFT_GRAPH[1080]};
					9'd185	:	PATTERN = {LEFT_GRAPH[1529], LEFT_GRAPH[1465], LEFT_GRAPH[1401], LEFT_GRAPH[1337], LEFT_GRAPH[1273], LEFT_GRAPH[1209], LEFT_GRAPH[1145], LEFT_GRAPH[1081]};
					9'd186	:	PATTERN = {LEFT_GRAPH[1530], LEFT_GRAPH[1466], LEFT_GRAPH[1402], LEFT_GRAPH[1338], LEFT_GRAPH[1274], LEFT_GRAPH[1210], LEFT_GRAPH[1146], LEFT_GRAPH[1082]};
					9'd187	:	PATTERN = {LEFT_GRAPH[1531], LEFT_GRAPH[1467], LEFT_GRAPH[1403], LEFT_GRAPH[1339], LEFT_GRAPH[1275], LEFT_GRAPH[1211], LEFT_GRAPH[1147], LEFT_GRAPH[1083]};
					9'd188	:	PATTERN = {LEFT_GRAPH[1532], LEFT_GRAPH[1468], LEFT_GRAPH[1404], LEFT_GRAPH[1340], LEFT_GRAPH[1276], LEFT_GRAPH[1212], LEFT_GRAPH[1148], LEFT_GRAPH[1084]};
					9'd189	:	PATTERN = {LEFT_GRAPH[1533], LEFT_GRAPH[1469], LEFT_GRAPH[1405], LEFT_GRAPH[1341], LEFT_GRAPH[1277], LEFT_GRAPH[1213], LEFT_GRAPH[1149], LEFT_GRAPH[1085]};
					9'd190	:	PATTERN = {LEFT_GRAPH[1534], LEFT_GRAPH[1470], LEFT_GRAPH[1406], LEFT_GRAPH[1342], LEFT_GRAPH[1278], LEFT_GRAPH[1214], LEFT_GRAPH[1150], LEFT_GRAPH[1086]};
					9'd191	:	PATTERN = {LEFT_GRAPH[1535], LEFT_GRAPH[1471], LEFT_GRAPH[1407], LEFT_GRAPH[1343], LEFT_GRAPH[1279], LEFT_GRAPH[1215], LEFT_GRAPH[1151], LEFT_GRAPH[1087]};
					9'd192	:	PATTERN = {LEFT_GRAPH[1984], LEFT_GRAPH[1920], LEFT_GRAPH[1856], LEFT_GRAPH[1792], LEFT_GRAPH[1728], LEFT_GRAPH[1664], LEFT_GRAPH[1600], LEFT_GRAPH[1536]};
					9'd193	:	PATTERN = {LEFT_GRAPH[1985], LEFT_GRAPH[1921], LEFT_GRAPH[1857], LEFT_GRAPH[1793], LEFT_GRAPH[1729], LEFT_GRAPH[1665], LEFT_GRAPH[1601], LEFT_GRAPH[1537]};
					9'd194	:	PATTERN = {LEFT_GRAPH[1986], LEFT_GRAPH[1922], LEFT_GRAPH[1858], LEFT_GRAPH[1794], LEFT_GRAPH[1730], LEFT_GRAPH[1666], LEFT_GRAPH[1602], LEFT_GRAPH[1538]};
					9'd195	:	PATTERN = {LEFT_GRAPH[1987], LEFT_GRAPH[1923], LEFT_GRAPH[1859], LEFT_GRAPH[1795], LEFT_GRAPH[1731], LEFT_GRAPH[1667], LEFT_GRAPH[1603], LEFT_GRAPH[1539]};
					9'd196	:	PATTERN = {LEFT_GRAPH[1988], LEFT_GRAPH[1924], LEFT_GRAPH[1860], LEFT_GRAPH[1796], LEFT_GRAPH[1732], LEFT_GRAPH[1668], LEFT_GRAPH[1604], LEFT_GRAPH[1540]};
					9'd197	:	PATTERN = {LEFT_GRAPH[1989], LEFT_GRAPH[1925], LEFT_GRAPH[1861], LEFT_GRAPH[1797], LEFT_GRAPH[1733], LEFT_GRAPH[1669], LEFT_GRAPH[1605], LEFT_GRAPH[1541]};
					9'd198	:	PATTERN = {LEFT_GRAPH[1990], LEFT_GRAPH[1926], LEFT_GRAPH[1862], LEFT_GRAPH[1798], LEFT_GRAPH[1734], LEFT_GRAPH[1670], LEFT_GRAPH[1606], LEFT_GRAPH[1542]};
					9'd199	:	PATTERN = {LEFT_GRAPH[1991], LEFT_GRAPH[1927], LEFT_GRAPH[1863], LEFT_GRAPH[1799], LEFT_GRAPH[1735], LEFT_GRAPH[1671], LEFT_GRAPH[1607], LEFT_GRAPH[1543]};
					9'd200	:	PATTERN = {LEFT_GRAPH[1992], LEFT_GRAPH[1928], LEFT_GRAPH[1864], LEFT_GRAPH[1800], LEFT_GRAPH[1736], LEFT_GRAPH[1672], LEFT_GRAPH[1608], LEFT_GRAPH[1544]};
					9'd201	:	PATTERN = {LEFT_GRAPH[1993], LEFT_GRAPH[1929], LEFT_GRAPH[1865], LEFT_GRAPH[1801], LEFT_GRAPH[1737], LEFT_GRAPH[1673], LEFT_GRAPH[1609], LEFT_GRAPH[1545]};
					9'd202	:	PATTERN = {LEFT_GRAPH[1994], LEFT_GRAPH[1930], LEFT_GRAPH[1866], LEFT_GRAPH[1802], LEFT_GRAPH[1738], LEFT_GRAPH[1674], LEFT_GRAPH[1610], LEFT_GRAPH[1546]};
					9'd203	:	PATTERN = {LEFT_GRAPH[1995], LEFT_GRAPH[1931], LEFT_GRAPH[1867], LEFT_GRAPH[1803], LEFT_GRAPH[1739], LEFT_GRAPH[1675], LEFT_GRAPH[1611], LEFT_GRAPH[1547]};
					9'd204	:	PATTERN = {LEFT_GRAPH[1996], LEFT_GRAPH[1932], LEFT_GRAPH[1868], LEFT_GRAPH[1804], LEFT_GRAPH[1740], LEFT_GRAPH[1676], LEFT_GRAPH[1612], LEFT_GRAPH[1548]};
					9'd205	:	PATTERN = {LEFT_GRAPH[1997], LEFT_GRAPH[1933], LEFT_GRAPH[1869], LEFT_GRAPH[1805], LEFT_GRAPH[1741], LEFT_GRAPH[1677], LEFT_GRAPH[1613], LEFT_GRAPH[1549]};
					9'd206	:	PATTERN = {LEFT_GRAPH[1998], LEFT_GRAPH[1934], LEFT_GRAPH[1870], LEFT_GRAPH[1806], LEFT_GRAPH[1742], LEFT_GRAPH[1678], LEFT_GRAPH[1614], LEFT_GRAPH[1550]};
					9'd207	:	PATTERN = {LEFT_GRAPH[1999], LEFT_GRAPH[1935], LEFT_GRAPH[1871], LEFT_GRAPH[1807], LEFT_GRAPH[1743], LEFT_GRAPH[1679], LEFT_GRAPH[1615], LEFT_GRAPH[1551]};
					9'd208	:	PATTERN = {LEFT_GRAPH[2000], LEFT_GRAPH[1936], LEFT_GRAPH[1872], LEFT_GRAPH[1808], LEFT_GRAPH[1744], LEFT_GRAPH[1680], LEFT_GRAPH[1616], LEFT_GRAPH[1552]};
					9'd209	:	PATTERN = {LEFT_GRAPH[2001], LEFT_GRAPH[1937], LEFT_GRAPH[1873], LEFT_GRAPH[1809], LEFT_GRAPH[1745], LEFT_GRAPH[1681], LEFT_GRAPH[1617], LEFT_GRAPH[1553]};
					9'd210	:	PATTERN = {LEFT_GRAPH[2002], LEFT_GRAPH[1938], LEFT_GRAPH[1874], LEFT_GRAPH[1810], LEFT_GRAPH[1746], LEFT_GRAPH[1682], LEFT_GRAPH[1618], LEFT_GRAPH[1554]};
					9'd211	:	PATTERN = {LEFT_GRAPH[2003], LEFT_GRAPH[1939], LEFT_GRAPH[1875], LEFT_GRAPH[1811], LEFT_GRAPH[1747], LEFT_GRAPH[1683], LEFT_GRAPH[1619], LEFT_GRAPH[1555]};
					9'd212	:	PATTERN = {LEFT_GRAPH[2004], LEFT_GRAPH[1940], LEFT_GRAPH[1876], LEFT_GRAPH[1812], LEFT_GRAPH[1748], LEFT_GRAPH[1684], LEFT_GRAPH[1620], LEFT_GRAPH[1556]};
					9'd213	:	PATTERN = {LEFT_GRAPH[2005], LEFT_GRAPH[1941], LEFT_GRAPH[1877], LEFT_GRAPH[1813], LEFT_GRAPH[1749], LEFT_GRAPH[1685], LEFT_GRAPH[1621], LEFT_GRAPH[1557]};
					9'd214	:	PATTERN = {LEFT_GRAPH[2006], LEFT_GRAPH[1942], LEFT_GRAPH[1878], LEFT_GRAPH[1814], LEFT_GRAPH[1750], LEFT_GRAPH[1686], LEFT_GRAPH[1622], LEFT_GRAPH[1558]};
					9'd215	:	PATTERN = {LEFT_GRAPH[2007], LEFT_GRAPH[1943], LEFT_GRAPH[1879], LEFT_GRAPH[1815], LEFT_GRAPH[1751], LEFT_GRAPH[1687], LEFT_GRAPH[1623], LEFT_GRAPH[1559]};
					9'd216	:	PATTERN = {LEFT_GRAPH[2008], LEFT_GRAPH[1944], LEFT_GRAPH[1880], LEFT_GRAPH[1816], LEFT_GRAPH[1752], LEFT_GRAPH[1688], LEFT_GRAPH[1624], LEFT_GRAPH[1560]};
					9'd217	:	PATTERN = {LEFT_GRAPH[2009], LEFT_GRAPH[1945], LEFT_GRAPH[1881], LEFT_GRAPH[1817], LEFT_GRAPH[1753], LEFT_GRAPH[1689], LEFT_GRAPH[1625], LEFT_GRAPH[1561]};
					9'd218	:	PATTERN = {LEFT_GRAPH[2010], LEFT_GRAPH[1946], LEFT_GRAPH[1882], LEFT_GRAPH[1818], LEFT_GRAPH[1754], LEFT_GRAPH[1690], LEFT_GRAPH[1626], LEFT_GRAPH[1562]};
					9'd219	:	PATTERN = {LEFT_GRAPH[2011], LEFT_GRAPH[1947], LEFT_GRAPH[1883], LEFT_GRAPH[1819], LEFT_GRAPH[1755], LEFT_GRAPH[1691], LEFT_GRAPH[1627], LEFT_GRAPH[1563]};
					9'd220	:	PATTERN = {LEFT_GRAPH[2012], LEFT_GRAPH[1948], LEFT_GRAPH[1884], LEFT_GRAPH[1820], LEFT_GRAPH[1756], LEFT_GRAPH[1692], LEFT_GRAPH[1628], LEFT_GRAPH[1564]};
					9'd221	:	PATTERN = {LEFT_GRAPH[2013], LEFT_GRAPH[1949], LEFT_GRAPH[1885], LEFT_GRAPH[1821], LEFT_GRAPH[1757], LEFT_GRAPH[1693], LEFT_GRAPH[1629], LEFT_GRAPH[1565]};
					9'd222	:	PATTERN = {LEFT_GRAPH[2014], LEFT_GRAPH[1950], LEFT_GRAPH[1886], LEFT_GRAPH[1822], LEFT_GRAPH[1758], LEFT_GRAPH[1694], LEFT_GRAPH[1630], LEFT_GRAPH[1566]};
					9'd223	:	PATTERN = {LEFT_GRAPH[2015], LEFT_GRAPH[1951], LEFT_GRAPH[1887], LEFT_GRAPH[1823], LEFT_GRAPH[1759], LEFT_GRAPH[1695], LEFT_GRAPH[1631], LEFT_GRAPH[1567]};
					9'd224	:	PATTERN = {LEFT_GRAPH[2016], LEFT_GRAPH[1952], LEFT_GRAPH[1888], LEFT_GRAPH[1824], LEFT_GRAPH[1760], LEFT_GRAPH[1696], LEFT_GRAPH[1632], LEFT_GRAPH[1568]};
					9'd225	:	PATTERN = {LEFT_GRAPH[2017], LEFT_GRAPH[1953], LEFT_GRAPH[1889], LEFT_GRAPH[1825], LEFT_GRAPH[1761], LEFT_GRAPH[1697], LEFT_GRAPH[1633], LEFT_GRAPH[1569]};
					9'd226	:	PATTERN = {LEFT_GRAPH[2018], LEFT_GRAPH[1954], LEFT_GRAPH[1890], LEFT_GRAPH[1826], LEFT_GRAPH[1762], LEFT_GRAPH[1698], LEFT_GRAPH[1634], LEFT_GRAPH[1570]};
					9'd227	:	PATTERN = {LEFT_GRAPH[2019], LEFT_GRAPH[1955], LEFT_GRAPH[1891], LEFT_GRAPH[1827], LEFT_GRAPH[1763], LEFT_GRAPH[1699], LEFT_GRAPH[1635], LEFT_GRAPH[1571]};
					9'd228	:	PATTERN = {LEFT_GRAPH[2020], LEFT_GRAPH[1956], LEFT_GRAPH[1892], LEFT_GRAPH[1828], LEFT_GRAPH[1764], LEFT_GRAPH[1700], LEFT_GRAPH[1636], LEFT_GRAPH[1572]};
					9'd229	:	PATTERN = {LEFT_GRAPH[2021], LEFT_GRAPH[1957], LEFT_GRAPH[1893], LEFT_GRAPH[1829], LEFT_GRAPH[1765], LEFT_GRAPH[1701], LEFT_GRAPH[1637], LEFT_GRAPH[1573]};
					9'd230	:	PATTERN = {LEFT_GRAPH[2022], LEFT_GRAPH[1958], LEFT_GRAPH[1894], LEFT_GRAPH[1830], LEFT_GRAPH[1766], LEFT_GRAPH[1702], LEFT_GRAPH[1638], LEFT_GRAPH[1574]};
					9'd231	:	PATTERN = {LEFT_GRAPH[2023], LEFT_GRAPH[1959], LEFT_GRAPH[1895], LEFT_GRAPH[1831], LEFT_GRAPH[1767], LEFT_GRAPH[1703], LEFT_GRAPH[1639], LEFT_GRAPH[1575]};
					9'd232	:	PATTERN = {LEFT_GRAPH[2024], LEFT_GRAPH[1960], LEFT_GRAPH[1896], LEFT_GRAPH[1832], LEFT_GRAPH[1768], LEFT_GRAPH[1704], LEFT_GRAPH[1640], LEFT_GRAPH[1576]};
					9'd233	:	PATTERN = {LEFT_GRAPH[2025], LEFT_GRAPH[1961], LEFT_GRAPH[1897], LEFT_GRAPH[1833], LEFT_GRAPH[1769], LEFT_GRAPH[1705], LEFT_GRAPH[1641], LEFT_GRAPH[1577]};
					9'd234	:	PATTERN = {LEFT_GRAPH[2026], LEFT_GRAPH[1962], LEFT_GRAPH[1898], LEFT_GRAPH[1834], LEFT_GRAPH[1770], LEFT_GRAPH[1706], LEFT_GRAPH[1642], LEFT_GRAPH[1578]};
					9'd235	:	PATTERN = {LEFT_GRAPH[2027], LEFT_GRAPH[1963], LEFT_GRAPH[1899], LEFT_GRAPH[1835], LEFT_GRAPH[1771], LEFT_GRAPH[1707], LEFT_GRAPH[1643], LEFT_GRAPH[1579]};
					9'd236	:	PATTERN = {LEFT_GRAPH[2028], LEFT_GRAPH[1964], LEFT_GRAPH[1900], LEFT_GRAPH[1836], LEFT_GRAPH[1772], LEFT_GRAPH[1708], LEFT_GRAPH[1644], LEFT_GRAPH[1580]};
					9'd237	:	PATTERN = {LEFT_GRAPH[2029], LEFT_GRAPH[1965], LEFT_GRAPH[1901], LEFT_GRAPH[1837], LEFT_GRAPH[1773], LEFT_GRAPH[1709], LEFT_GRAPH[1645], LEFT_GRAPH[1581]};
					9'd238	:	PATTERN = {LEFT_GRAPH[2030], LEFT_GRAPH[1966], LEFT_GRAPH[1902], LEFT_GRAPH[1838], LEFT_GRAPH[1774], LEFT_GRAPH[1710], LEFT_GRAPH[1646], LEFT_GRAPH[1582]};
					9'd239	:	PATTERN = {LEFT_GRAPH[2031], LEFT_GRAPH[1967], LEFT_GRAPH[1903], LEFT_GRAPH[1839], LEFT_GRAPH[1775], LEFT_GRAPH[1711], LEFT_GRAPH[1647], LEFT_GRAPH[1583]};
					9'd240	:	PATTERN = {LEFT_GRAPH[2032], LEFT_GRAPH[1968], LEFT_GRAPH[1904], LEFT_GRAPH[1840], LEFT_GRAPH[1776], LEFT_GRAPH[1712], LEFT_GRAPH[1648], LEFT_GRAPH[1584]};
					9'd241	:	PATTERN = {LEFT_GRAPH[2033], LEFT_GRAPH[1969], LEFT_GRAPH[1905], LEFT_GRAPH[1841], LEFT_GRAPH[1777], LEFT_GRAPH[1713], LEFT_GRAPH[1649], LEFT_GRAPH[1585]};
					9'd242	:	PATTERN = {LEFT_GRAPH[2034], LEFT_GRAPH[1970], LEFT_GRAPH[1906], LEFT_GRAPH[1842], LEFT_GRAPH[1778], LEFT_GRAPH[1714], LEFT_GRAPH[1650], LEFT_GRAPH[1586]};
					9'd243	:	PATTERN = {LEFT_GRAPH[2035], LEFT_GRAPH[1971], LEFT_GRAPH[1907], LEFT_GRAPH[1843], LEFT_GRAPH[1779], LEFT_GRAPH[1715], LEFT_GRAPH[1651], LEFT_GRAPH[1587]};
					9'd244	:	PATTERN = {LEFT_GRAPH[2036], LEFT_GRAPH[1972], LEFT_GRAPH[1908], LEFT_GRAPH[1844], LEFT_GRAPH[1780], LEFT_GRAPH[1716], LEFT_GRAPH[1652], LEFT_GRAPH[1588]};
					9'd245	:	PATTERN = {LEFT_GRAPH[2037], LEFT_GRAPH[1973], LEFT_GRAPH[1909], LEFT_GRAPH[1845], LEFT_GRAPH[1781], LEFT_GRAPH[1717], LEFT_GRAPH[1653], LEFT_GRAPH[1589]};
					9'd246	:	PATTERN = {LEFT_GRAPH[2038], LEFT_GRAPH[1974], LEFT_GRAPH[1910], LEFT_GRAPH[1846], LEFT_GRAPH[1782], LEFT_GRAPH[1718], LEFT_GRAPH[1654], LEFT_GRAPH[1590]};
					9'd247	:	PATTERN = {LEFT_GRAPH[2039], LEFT_GRAPH[1975], LEFT_GRAPH[1911], LEFT_GRAPH[1847], LEFT_GRAPH[1783], LEFT_GRAPH[1719], LEFT_GRAPH[1655], LEFT_GRAPH[1591]};
					9'd248	:	PATTERN = {LEFT_GRAPH[2040], LEFT_GRAPH[1976], LEFT_GRAPH[1912], LEFT_GRAPH[1848], LEFT_GRAPH[1784], LEFT_GRAPH[1720], LEFT_GRAPH[1656], LEFT_GRAPH[1592]};
					9'd249	:	PATTERN = {LEFT_GRAPH[2041], LEFT_GRAPH[1977], LEFT_GRAPH[1913], LEFT_GRAPH[1849], LEFT_GRAPH[1785], LEFT_GRAPH[1721], LEFT_GRAPH[1657], LEFT_GRAPH[1593]};
					9'd250	:	PATTERN = {LEFT_GRAPH[2042], LEFT_GRAPH[1978], LEFT_GRAPH[1914], LEFT_GRAPH[1850], LEFT_GRAPH[1786], LEFT_GRAPH[1722], LEFT_GRAPH[1658], LEFT_GRAPH[1594]};
					9'd251	:	PATTERN = {LEFT_GRAPH[2043], LEFT_GRAPH[1979], LEFT_GRAPH[1915], LEFT_GRAPH[1851], LEFT_GRAPH[1787], LEFT_GRAPH[1723], LEFT_GRAPH[1659], LEFT_GRAPH[1595]};
					9'd252	:	PATTERN = {LEFT_GRAPH[2044], LEFT_GRAPH[1980], LEFT_GRAPH[1916], LEFT_GRAPH[1852], LEFT_GRAPH[1788], LEFT_GRAPH[1724], LEFT_GRAPH[1660], LEFT_GRAPH[1596]};
					9'd253	:	PATTERN = {LEFT_GRAPH[2045], LEFT_GRAPH[1981], LEFT_GRAPH[1917], LEFT_GRAPH[1853], LEFT_GRAPH[1789], LEFT_GRAPH[1725], LEFT_GRAPH[1661], LEFT_GRAPH[1597]};
					9'd254	:	PATTERN = {LEFT_GRAPH[2046], LEFT_GRAPH[1982], LEFT_GRAPH[1918], LEFT_GRAPH[1854], LEFT_GRAPH[1790], LEFT_GRAPH[1726], LEFT_GRAPH[1662], LEFT_GRAPH[1598]};
					9'd255	:	PATTERN = {LEFT_GRAPH[2047], LEFT_GRAPH[1983], LEFT_GRAPH[1919], LEFT_GRAPH[1855], LEFT_GRAPH[1791], LEFT_GRAPH[1727], LEFT_GRAPH[1663], LEFT_GRAPH[1599]};
					9'd256	:	PATTERN = {LEFT_GRAPH[2496], LEFT_GRAPH[2432], LEFT_GRAPH[2368], LEFT_GRAPH[2304], LEFT_GRAPH[2240], LEFT_GRAPH[2176], LEFT_GRAPH[2112], LEFT_GRAPH[2048]};
					9'd257	:	PATTERN = {LEFT_GRAPH[2497], LEFT_GRAPH[2433], LEFT_GRAPH[2369], LEFT_GRAPH[2305], LEFT_GRAPH[2241], LEFT_GRAPH[2177], LEFT_GRAPH[2113], LEFT_GRAPH[2049]};
					9'd258	:	PATTERN = {LEFT_GRAPH[2498], LEFT_GRAPH[2434], LEFT_GRAPH[2370], LEFT_GRAPH[2306], LEFT_GRAPH[2242], LEFT_GRAPH[2178], LEFT_GRAPH[2114], LEFT_GRAPH[2050]};
					9'd259	:	PATTERN = {LEFT_GRAPH[2499], LEFT_GRAPH[2435], LEFT_GRAPH[2371], LEFT_GRAPH[2307], LEFT_GRAPH[2243], LEFT_GRAPH[2179], LEFT_GRAPH[2115], LEFT_GRAPH[2051]};
					9'd260	:	PATTERN = {LEFT_GRAPH[2500], LEFT_GRAPH[2436], LEFT_GRAPH[2372], LEFT_GRAPH[2308], LEFT_GRAPH[2244], LEFT_GRAPH[2180], LEFT_GRAPH[2116], LEFT_GRAPH[2052]};
					9'd261	:	PATTERN = {LEFT_GRAPH[2501], LEFT_GRAPH[2437], LEFT_GRAPH[2373], LEFT_GRAPH[2309], LEFT_GRAPH[2245], LEFT_GRAPH[2181], LEFT_GRAPH[2117], LEFT_GRAPH[2053]};
					9'd262	:	PATTERN = {LEFT_GRAPH[2502], LEFT_GRAPH[2438], LEFT_GRAPH[2374], LEFT_GRAPH[2310], LEFT_GRAPH[2246], LEFT_GRAPH[2182], LEFT_GRAPH[2118], LEFT_GRAPH[2054]};
					9'd263	:	PATTERN = {LEFT_GRAPH[2503], LEFT_GRAPH[2439], LEFT_GRAPH[2375], LEFT_GRAPH[2311], LEFT_GRAPH[2247], LEFT_GRAPH[2183], LEFT_GRAPH[2119], LEFT_GRAPH[2055]};
					9'd264	:	PATTERN = {LEFT_GRAPH[2504], LEFT_GRAPH[2440], LEFT_GRAPH[2376], LEFT_GRAPH[2312], LEFT_GRAPH[2248], LEFT_GRAPH[2184], LEFT_GRAPH[2120], LEFT_GRAPH[2056]};
					9'd265	:	PATTERN = {LEFT_GRAPH[2505], LEFT_GRAPH[2441], LEFT_GRAPH[2377], LEFT_GRAPH[2313], LEFT_GRAPH[2249], LEFT_GRAPH[2185], LEFT_GRAPH[2121], LEFT_GRAPH[2057]};
					9'd266	:	PATTERN = {LEFT_GRAPH[2506], LEFT_GRAPH[2442], LEFT_GRAPH[2378], LEFT_GRAPH[2314], LEFT_GRAPH[2250], LEFT_GRAPH[2186], LEFT_GRAPH[2122], LEFT_GRAPH[2058]};
					9'd267	:	PATTERN = {LEFT_GRAPH[2507], LEFT_GRAPH[2443], LEFT_GRAPH[2379], LEFT_GRAPH[2315], LEFT_GRAPH[2251], LEFT_GRAPH[2187], LEFT_GRAPH[2123], LEFT_GRAPH[2059]};
					9'd268	:	PATTERN = {LEFT_GRAPH[2508], LEFT_GRAPH[2444], LEFT_GRAPH[2380], LEFT_GRAPH[2316], LEFT_GRAPH[2252], LEFT_GRAPH[2188], LEFT_GRAPH[2124], LEFT_GRAPH[2060]};
					9'd269	:	PATTERN = {LEFT_GRAPH[2509], LEFT_GRAPH[2445], LEFT_GRAPH[2381], LEFT_GRAPH[2317], LEFT_GRAPH[2253], LEFT_GRAPH[2189], LEFT_GRAPH[2125], LEFT_GRAPH[2061]};
					9'd270	:	PATTERN = {LEFT_GRAPH[2510], LEFT_GRAPH[2446], LEFT_GRAPH[2382], LEFT_GRAPH[2318], LEFT_GRAPH[2254], LEFT_GRAPH[2190], LEFT_GRAPH[2126], LEFT_GRAPH[2062]};
					9'd271	:	PATTERN = {LEFT_GRAPH[2511], LEFT_GRAPH[2447], LEFT_GRAPH[2383], LEFT_GRAPH[2319], LEFT_GRAPH[2255], LEFT_GRAPH[2191], LEFT_GRAPH[2127], LEFT_GRAPH[2063]};
					9'd272	:	PATTERN = {LEFT_GRAPH[2512], LEFT_GRAPH[2448], LEFT_GRAPH[2384], LEFT_GRAPH[2320], LEFT_GRAPH[2256], LEFT_GRAPH[2192], LEFT_GRAPH[2128], LEFT_GRAPH[2064]};
					9'd273	:	PATTERN = {LEFT_GRAPH[2513], LEFT_GRAPH[2449], LEFT_GRAPH[2385], LEFT_GRAPH[2321], LEFT_GRAPH[2257], LEFT_GRAPH[2193], LEFT_GRAPH[2129], LEFT_GRAPH[2065]};
					9'd274	:	PATTERN = {LEFT_GRAPH[2514], LEFT_GRAPH[2450], LEFT_GRAPH[2386], LEFT_GRAPH[2322], LEFT_GRAPH[2258], LEFT_GRAPH[2194], LEFT_GRAPH[2130], LEFT_GRAPH[2066]};
					9'd275	:	PATTERN = {LEFT_GRAPH[2515], LEFT_GRAPH[2451], LEFT_GRAPH[2387], LEFT_GRAPH[2323], LEFT_GRAPH[2259], LEFT_GRAPH[2195], LEFT_GRAPH[2131], LEFT_GRAPH[2067]};
					9'd276	:	PATTERN = {LEFT_GRAPH[2516], LEFT_GRAPH[2452], LEFT_GRAPH[2388], LEFT_GRAPH[2324], LEFT_GRAPH[2260], LEFT_GRAPH[2196], LEFT_GRAPH[2132], LEFT_GRAPH[2068]};
					9'd277	:	PATTERN = {LEFT_GRAPH[2517], LEFT_GRAPH[2453], LEFT_GRAPH[2389], LEFT_GRAPH[2325], LEFT_GRAPH[2261], LEFT_GRAPH[2197], LEFT_GRAPH[2133], LEFT_GRAPH[2069]};
					9'd278	:	PATTERN = {LEFT_GRAPH[2518], LEFT_GRAPH[2454], LEFT_GRAPH[2390], LEFT_GRAPH[2326], LEFT_GRAPH[2262], LEFT_GRAPH[2198], LEFT_GRAPH[2134], LEFT_GRAPH[2070]};
					9'd279	:	PATTERN = {LEFT_GRAPH[2519], LEFT_GRAPH[2455], LEFT_GRAPH[2391], LEFT_GRAPH[2327], LEFT_GRAPH[2263], LEFT_GRAPH[2199], LEFT_GRAPH[2135], LEFT_GRAPH[2071]};
					9'd280	:	PATTERN = {LEFT_GRAPH[2520], LEFT_GRAPH[2456], LEFT_GRAPH[2392], LEFT_GRAPH[2328], LEFT_GRAPH[2264], LEFT_GRAPH[2200], LEFT_GRAPH[2136], LEFT_GRAPH[2072]};
					9'd281	:	PATTERN = {LEFT_GRAPH[2521], LEFT_GRAPH[2457], LEFT_GRAPH[2393], LEFT_GRAPH[2329], LEFT_GRAPH[2265], LEFT_GRAPH[2201], LEFT_GRAPH[2137], LEFT_GRAPH[2073]};
					9'd282	:	PATTERN = {LEFT_GRAPH[2522], LEFT_GRAPH[2458], LEFT_GRAPH[2394], LEFT_GRAPH[2330], LEFT_GRAPH[2266], LEFT_GRAPH[2202], LEFT_GRAPH[2138], LEFT_GRAPH[2074]};
					9'd283	:	PATTERN = {LEFT_GRAPH[2523], LEFT_GRAPH[2459], LEFT_GRAPH[2395], LEFT_GRAPH[2331], LEFT_GRAPH[2267], LEFT_GRAPH[2203], LEFT_GRAPH[2139], LEFT_GRAPH[2075]};
					9'd284	:	PATTERN = {LEFT_GRAPH[2524], LEFT_GRAPH[2460], LEFT_GRAPH[2396], LEFT_GRAPH[2332], LEFT_GRAPH[2268], LEFT_GRAPH[2204], LEFT_GRAPH[2140], LEFT_GRAPH[2076]};
					9'd285	:	PATTERN = {LEFT_GRAPH[2525], LEFT_GRAPH[2461], LEFT_GRAPH[2397], LEFT_GRAPH[2333], LEFT_GRAPH[2269], LEFT_GRAPH[2205], LEFT_GRAPH[2141], LEFT_GRAPH[2077]};
					9'd286	:	PATTERN = {LEFT_GRAPH[2526], LEFT_GRAPH[2462], LEFT_GRAPH[2398], LEFT_GRAPH[2334], LEFT_GRAPH[2270], LEFT_GRAPH[2206], LEFT_GRAPH[2142], LEFT_GRAPH[2078]};
					9'd287	:	PATTERN = {LEFT_GRAPH[2527], LEFT_GRAPH[2463], LEFT_GRAPH[2399], LEFT_GRAPH[2335], LEFT_GRAPH[2271], LEFT_GRAPH[2207], LEFT_GRAPH[2143], LEFT_GRAPH[2079]};
					9'd288	:	PATTERN = {LEFT_GRAPH[2528], LEFT_GRAPH[2464], LEFT_GRAPH[2400], LEFT_GRAPH[2336], LEFT_GRAPH[2272], LEFT_GRAPH[2208], LEFT_GRAPH[2144], LEFT_GRAPH[2080]};
					9'd289	:	PATTERN = {LEFT_GRAPH[2529], LEFT_GRAPH[2465], LEFT_GRAPH[2401], LEFT_GRAPH[2337], LEFT_GRAPH[2273], LEFT_GRAPH[2209], LEFT_GRAPH[2145], LEFT_GRAPH[2081]};
					9'd290	:	PATTERN = {LEFT_GRAPH[2530], LEFT_GRAPH[2466], LEFT_GRAPH[2402], LEFT_GRAPH[2338], LEFT_GRAPH[2274], LEFT_GRAPH[2210], LEFT_GRAPH[2146], LEFT_GRAPH[2082]};
					9'd291	:	PATTERN = {LEFT_GRAPH[2531], LEFT_GRAPH[2467], LEFT_GRAPH[2403], LEFT_GRAPH[2339], LEFT_GRAPH[2275], LEFT_GRAPH[2211], LEFT_GRAPH[2147], LEFT_GRAPH[2083]};
					9'd292	:	PATTERN = {LEFT_GRAPH[2532], LEFT_GRAPH[2468], LEFT_GRAPH[2404], LEFT_GRAPH[2340], LEFT_GRAPH[2276], LEFT_GRAPH[2212], LEFT_GRAPH[2148], LEFT_GRAPH[2084]};
					9'd293	:	PATTERN = {LEFT_GRAPH[2533], LEFT_GRAPH[2469], LEFT_GRAPH[2405], LEFT_GRAPH[2341], LEFT_GRAPH[2277], LEFT_GRAPH[2213], LEFT_GRAPH[2149], LEFT_GRAPH[2085]};
					9'd294	:	PATTERN = {LEFT_GRAPH[2534], LEFT_GRAPH[2470], LEFT_GRAPH[2406], LEFT_GRAPH[2342], LEFT_GRAPH[2278], LEFT_GRAPH[2214], LEFT_GRAPH[2150], LEFT_GRAPH[2086]};
					9'd295	:	PATTERN = {LEFT_GRAPH[2535], LEFT_GRAPH[2471], LEFT_GRAPH[2407], LEFT_GRAPH[2343], LEFT_GRAPH[2279], LEFT_GRAPH[2215], LEFT_GRAPH[2151], LEFT_GRAPH[2087]};
					9'd296	:	PATTERN = {LEFT_GRAPH[2536], LEFT_GRAPH[2472], LEFT_GRAPH[2408], LEFT_GRAPH[2344], LEFT_GRAPH[2280], LEFT_GRAPH[2216], LEFT_GRAPH[2152], LEFT_GRAPH[2088]};
					9'd297	:	PATTERN = {LEFT_GRAPH[2537], LEFT_GRAPH[2473], LEFT_GRAPH[2409], LEFT_GRAPH[2345], LEFT_GRAPH[2281], LEFT_GRAPH[2217], LEFT_GRAPH[2153], LEFT_GRAPH[2089]};
					9'd298	:	PATTERN = {LEFT_GRAPH[2538], LEFT_GRAPH[2474], LEFT_GRAPH[2410], LEFT_GRAPH[2346], LEFT_GRAPH[2282], LEFT_GRAPH[2218], LEFT_GRAPH[2154], LEFT_GRAPH[2090]};
					9'd299	:	PATTERN = {LEFT_GRAPH[2539], LEFT_GRAPH[2475], LEFT_GRAPH[2411], LEFT_GRAPH[2347], LEFT_GRAPH[2283], LEFT_GRAPH[2219], LEFT_GRAPH[2155], LEFT_GRAPH[2091]};
					9'd300	:	PATTERN = {LEFT_GRAPH[2540], LEFT_GRAPH[2476], LEFT_GRAPH[2412], LEFT_GRAPH[2348], LEFT_GRAPH[2284], LEFT_GRAPH[2220], LEFT_GRAPH[2156], LEFT_GRAPH[2092]};
					9'd301	:	PATTERN = {LEFT_GRAPH[2541], LEFT_GRAPH[2477], LEFT_GRAPH[2413], LEFT_GRAPH[2349], LEFT_GRAPH[2285], LEFT_GRAPH[2221], LEFT_GRAPH[2157], LEFT_GRAPH[2093]};
					9'd302	:	PATTERN = {LEFT_GRAPH[2542], LEFT_GRAPH[2478], LEFT_GRAPH[2414], LEFT_GRAPH[2350], LEFT_GRAPH[2286], LEFT_GRAPH[2222], LEFT_GRAPH[2158], LEFT_GRAPH[2094]};
					9'd303	:	PATTERN = {LEFT_GRAPH[2543], LEFT_GRAPH[2479], LEFT_GRAPH[2415], LEFT_GRAPH[2351], LEFT_GRAPH[2287], LEFT_GRAPH[2223], LEFT_GRAPH[2159], LEFT_GRAPH[2095]};
					9'd304	:	PATTERN = {LEFT_GRAPH[2544], LEFT_GRAPH[2480], LEFT_GRAPH[2416], LEFT_GRAPH[2352], LEFT_GRAPH[2288], LEFT_GRAPH[2224], LEFT_GRAPH[2160], LEFT_GRAPH[2096]};
					9'd305	:	PATTERN = {LEFT_GRAPH[2545], LEFT_GRAPH[2481], LEFT_GRAPH[2417], LEFT_GRAPH[2353], LEFT_GRAPH[2289], LEFT_GRAPH[2225], LEFT_GRAPH[2161], LEFT_GRAPH[2097]};
					9'd306	:	PATTERN = {LEFT_GRAPH[2546], LEFT_GRAPH[2482], LEFT_GRAPH[2418], LEFT_GRAPH[2354], LEFT_GRAPH[2290], LEFT_GRAPH[2226], LEFT_GRAPH[2162], LEFT_GRAPH[2098]};
					9'd307	:	PATTERN = {LEFT_GRAPH[2547], LEFT_GRAPH[2483], LEFT_GRAPH[2419], LEFT_GRAPH[2355], LEFT_GRAPH[2291], LEFT_GRAPH[2227], LEFT_GRAPH[2163], LEFT_GRAPH[2099]};
					9'd308	:	PATTERN = {LEFT_GRAPH[2548], LEFT_GRAPH[2484], LEFT_GRAPH[2420], LEFT_GRAPH[2356], LEFT_GRAPH[2292], LEFT_GRAPH[2228], LEFT_GRAPH[2164], LEFT_GRAPH[2100]};
					9'd309	:	PATTERN = {LEFT_GRAPH[2549], LEFT_GRAPH[2485], LEFT_GRAPH[2421], LEFT_GRAPH[2357], LEFT_GRAPH[2293], LEFT_GRAPH[2229], LEFT_GRAPH[2165], LEFT_GRAPH[2101]};
					9'd310	:	PATTERN = {LEFT_GRAPH[2550], LEFT_GRAPH[2486], LEFT_GRAPH[2422], LEFT_GRAPH[2358], LEFT_GRAPH[2294], LEFT_GRAPH[2230], LEFT_GRAPH[2166], LEFT_GRAPH[2102]};
					9'd311	:	PATTERN = {LEFT_GRAPH[2551], LEFT_GRAPH[2487], LEFT_GRAPH[2423], LEFT_GRAPH[2359], LEFT_GRAPH[2295], LEFT_GRAPH[2231], LEFT_GRAPH[2167], LEFT_GRAPH[2103]};
					9'd312	:	PATTERN = {LEFT_GRAPH[2552], LEFT_GRAPH[2488], LEFT_GRAPH[2424], LEFT_GRAPH[2360], LEFT_GRAPH[2296], LEFT_GRAPH[2232], LEFT_GRAPH[2168], LEFT_GRAPH[2104]};
					9'd313	:	PATTERN = {LEFT_GRAPH[2553], LEFT_GRAPH[2489], LEFT_GRAPH[2425], LEFT_GRAPH[2361], LEFT_GRAPH[2297], LEFT_GRAPH[2233], LEFT_GRAPH[2169], LEFT_GRAPH[2105]};
					9'd314	:	PATTERN = {LEFT_GRAPH[2554], LEFT_GRAPH[2490], LEFT_GRAPH[2426], LEFT_GRAPH[2362], LEFT_GRAPH[2298], LEFT_GRAPH[2234], LEFT_GRAPH[2170], LEFT_GRAPH[2106]};
					9'd315	:	PATTERN = {LEFT_GRAPH[2555], LEFT_GRAPH[2491], LEFT_GRAPH[2427], LEFT_GRAPH[2363], LEFT_GRAPH[2299], LEFT_GRAPH[2235], LEFT_GRAPH[2171], LEFT_GRAPH[2107]};
					9'd316	:	PATTERN = {LEFT_GRAPH[2556], LEFT_GRAPH[2492], LEFT_GRAPH[2428], LEFT_GRAPH[2364], LEFT_GRAPH[2300], LEFT_GRAPH[2236], LEFT_GRAPH[2172], LEFT_GRAPH[2108]};
					9'd317	:	PATTERN = {LEFT_GRAPH[2557], LEFT_GRAPH[2493], LEFT_GRAPH[2429], LEFT_GRAPH[2365], LEFT_GRAPH[2301], LEFT_GRAPH[2237], LEFT_GRAPH[2173], LEFT_GRAPH[2109]};
					9'd318	:	PATTERN = {LEFT_GRAPH[2558], LEFT_GRAPH[2494], LEFT_GRAPH[2430], LEFT_GRAPH[2366], LEFT_GRAPH[2302], LEFT_GRAPH[2238], LEFT_GRAPH[2174], LEFT_GRAPH[2110]};
					9'd319	:	PATTERN = {LEFT_GRAPH[2559], LEFT_GRAPH[2495], LEFT_GRAPH[2431], LEFT_GRAPH[2367], LEFT_GRAPH[2303], LEFT_GRAPH[2239], LEFT_GRAPH[2175], LEFT_GRAPH[2111]};
					9'd320	:	PATTERN = {LEFT_GRAPH[3008], LEFT_GRAPH[2944], LEFT_GRAPH[2880], LEFT_GRAPH[2816], LEFT_GRAPH[2752], LEFT_GRAPH[2688], LEFT_GRAPH[2624], LEFT_GRAPH[2560]};
					9'd321	:	PATTERN = {LEFT_GRAPH[3009], LEFT_GRAPH[2945], LEFT_GRAPH[2881], LEFT_GRAPH[2817], LEFT_GRAPH[2753], LEFT_GRAPH[2689], LEFT_GRAPH[2625], LEFT_GRAPH[2561]};
					9'd322	:	PATTERN = {LEFT_GRAPH[3010], LEFT_GRAPH[2946], LEFT_GRAPH[2882], LEFT_GRAPH[2818], LEFT_GRAPH[2754], LEFT_GRAPH[2690], LEFT_GRAPH[2626], LEFT_GRAPH[2562]};
					9'd323	:	PATTERN = {LEFT_GRAPH[3011], LEFT_GRAPH[2947], LEFT_GRAPH[2883], LEFT_GRAPH[2819], LEFT_GRAPH[2755], LEFT_GRAPH[2691], LEFT_GRAPH[2627], LEFT_GRAPH[2563]};
					9'd324	:	PATTERN = {LEFT_GRAPH[3012], LEFT_GRAPH[2948], LEFT_GRAPH[2884], LEFT_GRAPH[2820], LEFT_GRAPH[2756], LEFT_GRAPH[2692], LEFT_GRAPH[2628], LEFT_GRAPH[2564]};
					9'd325	:	PATTERN = {LEFT_GRAPH[3013], LEFT_GRAPH[2949], LEFT_GRAPH[2885], LEFT_GRAPH[2821], LEFT_GRAPH[2757], LEFT_GRAPH[2693], LEFT_GRAPH[2629], LEFT_GRAPH[2565]};
					9'd326	:	PATTERN = {LEFT_GRAPH[3014], LEFT_GRAPH[2950], LEFT_GRAPH[2886], LEFT_GRAPH[2822], LEFT_GRAPH[2758], LEFT_GRAPH[2694], LEFT_GRAPH[2630], LEFT_GRAPH[2566]};
					9'd327	:	PATTERN = {LEFT_GRAPH[3015], LEFT_GRAPH[2951], LEFT_GRAPH[2887], LEFT_GRAPH[2823], LEFT_GRAPH[2759], LEFT_GRAPH[2695], LEFT_GRAPH[2631], LEFT_GRAPH[2567]};
					9'd328	:	PATTERN = {LEFT_GRAPH[3016], LEFT_GRAPH[2952], LEFT_GRAPH[2888], LEFT_GRAPH[2824], LEFT_GRAPH[2760], LEFT_GRAPH[2696], LEFT_GRAPH[2632], LEFT_GRAPH[2568]};
					9'd329	:	PATTERN = {LEFT_GRAPH[3017], LEFT_GRAPH[2953], LEFT_GRAPH[2889], LEFT_GRAPH[2825], LEFT_GRAPH[2761], LEFT_GRAPH[2697], LEFT_GRAPH[2633], LEFT_GRAPH[2569]};
					9'd330	:	PATTERN = {LEFT_GRAPH[3018], LEFT_GRAPH[2954], LEFT_GRAPH[2890], LEFT_GRAPH[2826], LEFT_GRAPH[2762], LEFT_GRAPH[2698], LEFT_GRAPH[2634], LEFT_GRAPH[2570]};
					9'd331	:	PATTERN = {LEFT_GRAPH[3019], LEFT_GRAPH[2955], LEFT_GRAPH[2891], LEFT_GRAPH[2827], LEFT_GRAPH[2763], LEFT_GRAPH[2699], LEFT_GRAPH[2635], LEFT_GRAPH[2571]};
					9'd332	:	PATTERN = {LEFT_GRAPH[3020], LEFT_GRAPH[2956], LEFT_GRAPH[2892], LEFT_GRAPH[2828], LEFT_GRAPH[2764], LEFT_GRAPH[2700], LEFT_GRAPH[2636], LEFT_GRAPH[2572]};
					9'd333	:	PATTERN = {LEFT_GRAPH[3021], LEFT_GRAPH[2957], LEFT_GRAPH[2893], LEFT_GRAPH[2829], LEFT_GRAPH[2765], LEFT_GRAPH[2701], LEFT_GRAPH[2637], LEFT_GRAPH[2573]};
					9'd334	:	PATTERN = {LEFT_GRAPH[3022], LEFT_GRAPH[2958], LEFT_GRAPH[2894], LEFT_GRAPH[2830], LEFT_GRAPH[2766], LEFT_GRAPH[2702], LEFT_GRAPH[2638], LEFT_GRAPH[2574]};
					9'd335	:	PATTERN = {LEFT_GRAPH[3023], LEFT_GRAPH[2959], LEFT_GRAPH[2895], LEFT_GRAPH[2831], LEFT_GRAPH[2767], LEFT_GRAPH[2703], LEFT_GRAPH[2639], LEFT_GRAPH[2575]};
					9'd336	:	PATTERN = {LEFT_GRAPH[3024], LEFT_GRAPH[2960], LEFT_GRAPH[2896], LEFT_GRAPH[2832], LEFT_GRAPH[2768], LEFT_GRAPH[2704], LEFT_GRAPH[2640], LEFT_GRAPH[2576]};
					9'd337	:	PATTERN = {LEFT_GRAPH[3025], LEFT_GRAPH[2961], LEFT_GRAPH[2897], LEFT_GRAPH[2833], LEFT_GRAPH[2769], LEFT_GRAPH[2705], LEFT_GRAPH[2641], LEFT_GRAPH[2577]};
					9'd338	:	PATTERN = {LEFT_GRAPH[3026], LEFT_GRAPH[2962], LEFT_GRAPH[2898], LEFT_GRAPH[2834], LEFT_GRAPH[2770], LEFT_GRAPH[2706], LEFT_GRAPH[2642], LEFT_GRAPH[2578]};
					9'd339	:	PATTERN = {LEFT_GRAPH[3027], LEFT_GRAPH[2963], LEFT_GRAPH[2899], LEFT_GRAPH[2835], LEFT_GRAPH[2771], LEFT_GRAPH[2707], LEFT_GRAPH[2643], LEFT_GRAPH[2579]};
					9'd340	:	PATTERN = {LEFT_GRAPH[3028], LEFT_GRAPH[2964], LEFT_GRAPH[2900], LEFT_GRAPH[2836], LEFT_GRAPH[2772], LEFT_GRAPH[2708], LEFT_GRAPH[2644], LEFT_GRAPH[2580]};
					9'd341	:	PATTERN = {LEFT_GRAPH[3029], LEFT_GRAPH[2965], LEFT_GRAPH[2901], LEFT_GRAPH[2837], LEFT_GRAPH[2773], LEFT_GRAPH[2709], LEFT_GRAPH[2645], LEFT_GRAPH[2581]};
					9'd342	:	PATTERN = {LEFT_GRAPH[3030], LEFT_GRAPH[2966], LEFT_GRAPH[2902], LEFT_GRAPH[2838], LEFT_GRAPH[2774], LEFT_GRAPH[2710], LEFT_GRAPH[2646], LEFT_GRAPH[2582]};
					9'd343	:	PATTERN = {LEFT_GRAPH[3031], LEFT_GRAPH[2967], LEFT_GRAPH[2903], LEFT_GRAPH[2839], LEFT_GRAPH[2775], LEFT_GRAPH[2711], LEFT_GRAPH[2647], LEFT_GRAPH[2583]};
					9'd344	:	PATTERN = {LEFT_GRAPH[3032], LEFT_GRAPH[2968], LEFT_GRAPH[2904], LEFT_GRAPH[2840], LEFT_GRAPH[2776], LEFT_GRAPH[2712], LEFT_GRAPH[2648], LEFT_GRAPH[2584]};
					9'd345	:	PATTERN = {LEFT_GRAPH[3033], LEFT_GRAPH[2969], LEFT_GRAPH[2905], LEFT_GRAPH[2841], LEFT_GRAPH[2777], LEFT_GRAPH[2713], LEFT_GRAPH[2649], LEFT_GRAPH[2585]};
					9'd346	:	PATTERN = {LEFT_GRAPH[3034], LEFT_GRAPH[2970], LEFT_GRAPH[2906], LEFT_GRAPH[2842], LEFT_GRAPH[2778], LEFT_GRAPH[2714], LEFT_GRAPH[2650], LEFT_GRAPH[2586]};
					9'd347	:	PATTERN = {LEFT_GRAPH[3035], LEFT_GRAPH[2971], LEFT_GRAPH[2907], LEFT_GRAPH[2843], LEFT_GRAPH[2779], LEFT_GRAPH[2715], LEFT_GRAPH[2651], LEFT_GRAPH[2587]};
					9'd348	:	PATTERN = {LEFT_GRAPH[3036], LEFT_GRAPH[2972], LEFT_GRAPH[2908], LEFT_GRAPH[2844], LEFT_GRAPH[2780], LEFT_GRAPH[2716], LEFT_GRAPH[2652], LEFT_GRAPH[2588]};
					9'd349	:	PATTERN = {LEFT_GRAPH[3037], LEFT_GRAPH[2973], LEFT_GRAPH[2909], LEFT_GRAPH[2845], LEFT_GRAPH[2781], LEFT_GRAPH[2717], LEFT_GRAPH[2653], LEFT_GRAPH[2589]};
					9'd350	:	PATTERN = {LEFT_GRAPH[3038], LEFT_GRAPH[2974], LEFT_GRAPH[2910], LEFT_GRAPH[2846], LEFT_GRAPH[2782], LEFT_GRAPH[2718], LEFT_GRAPH[2654], LEFT_GRAPH[2590]};
					9'd351	:	PATTERN = {LEFT_GRAPH[3039], LEFT_GRAPH[2975], LEFT_GRAPH[2911], LEFT_GRAPH[2847], LEFT_GRAPH[2783], LEFT_GRAPH[2719], LEFT_GRAPH[2655], LEFT_GRAPH[2591]};
					9'd352	:	PATTERN = {LEFT_GRAPH[3040], LEFT_GRAPH[2976], LEFT_GRAPH[2912], LEFT_GRAPH[2848], LEFT_GRAPH[2784], LEFT_GRAPH[2720], LEFT_GRAPH[2656], LEFT_GRAPH[2592]};
					9'd353	:	PATTERN = {LEFT_GRAPH[3041], LEFT_GRAPH[2977], LEFT_GRAPH[2913], LEFT_GRAPH[2849], LEFT_GRAPH[2785], LEFT_GRAPH[2721], LEFT_GRAPH[2657], LEFT_GRAPH[2593]};
					9'd354	:	PATTERN = {LEFT_GRAPH[3042], LEFT_GRAPH[2978], LEFT_GRAPH[2914], LEFT_GRAPH[2850], LEFT_GRAPH[2786], LEFT_GRAPH[2722], LEFT_GRAPH[2658], LEFT_GRAPH[2594]};
					9'd355	:	PATTERN = {LEFT_GRAPH[3043], LEFT_GRAPH[2979], LEFT_GRAPH[2915], LEFT_GRAPH[2851], LEFT_GRAPH[2787], LEFT_GRAPH[2723], LEFT_GRAPH[2659], LEFT_GRAPH[2595]};
					9'd356	:	PATTERN = {LEFT_GRAPH[3044], LEFT_GRAPH[2980], LEFT_GRAPH[2916], LEFT_GRAPH[2852], LEFT_GRAPH[2788], LEFT_GRAPH[2724], LEFT_GRAPH[2660], LEFT_GRAPH[2596]};
					9'd357	:	PATTERN = {LEFT_GRAPH[3045], LEFT_GRAPH[2981], LEFT_GRAPH[2917], LEFT_GRAPH[2853], LEFT_GRAPH[2789], LEFT_GRAPH[2725], LEFT_GRAPH[2661], LEFT_GRAPH[2597]};
					9'd358	:	PATTERN = {LEFT_GRAPH[3046], LEFT_GRAPH[2982], LEFT_GRAPH[2918], LEFT_GRAPH[2854], LEFT_GRAPH[2790], LEFT_GRAPH[2726], LEFT_GRAPH[2662], LEFT_GRAPH[2598]};
					9'd359	:	PATTERN = {LEFT_GRAPH[3047], LEFT_GRAPH[2983], LEFT_GRAPH[2919], LEFT_GRAPH[2855], LEFT_GRAPH[2791], LEFT_GRAPH[2727], LEFT_GRAPH[2663], LEFT_GRAPH[2599]};
					9'd360	:	PATTERN = {LEFT_GRAPH[3048], LEFT_GRAPH[2984], LEFT_GRAPH[2920], LEFT_GRAPH[2856], LEFT_GRAPH[2792], LEFT_GRAPH[2728], LEFT_GRAPH[2664], LEFT_GRAPH[2600]};
					9'd361	:	PATTERN = {LEFT_GRAPH[3049], LEFT_GRAPH[2985], LEFT_GRAPH[2921], LEFT_GRAPH[2857], LEFT_GRAPH[2793], LEFT_GRAPH[2729], LEFT_GRAPH[2665], LEFT_GRAPH[2601]};
					9'd362	:	PATTERN = {LEFT_GRAPH[3050], LEFT_GRAPH[2986], LEFT_GRAPH[2922], LEFT_GRAPH[2858], LEFT_GRAPH[2794], LEFT_GRAPH[2730], LEFT_GRAPH[2666], LEFT_GRAPH[2602]};
					9'd363	:	PATTERN = {LEFT_GRAPH[3051], LEFT_GRAPH[2987], LEFT_GRAPH[2923], LEFT_GRAPH[2859], LEFT_GRAPH[2795], LEFT_GRAPH[2731], LEFT_GRAPH[2667], LEFT_GRAPH[2603]};
					9'd364	:	PATTERN = {LEFT_GRAPH[3052], LEFT_GRAPH[2988], LEFT_GRAPH[2924], LEFT_GRAPH[2860], LEFT_GRAPH[2796], LEFT_GRAPH[2732], LEFT_GRAPH[2668], LEFT_GRAPH[2604]};
					9'd365	:	PATTERN = {LEFT_GRAPH[3053], LEFT_GRAPH[2989], LEFT_GRAPH[2925], LEFT_GRAPH[2861], LEFT_GRAPH[2797], LEFT_GRAPH[2733], LEFT_GRAPH[2669], LEFT_GRAPH[2605]};
					9'd366	:	PATTERN = {LEFT_GRAPH[3054], LEFT_GRAPH[2990], LEFT_GRAPH[2926], LEFT_GRAPH[2862], LEFT_GRAPH[2798], LEFT_GRAPH[2734], LEFT_GRAPH[2670], LEFT_GRAPH[2606]};
					9'd367	:	PATTERN = {LEFT_GRAPH[3055], LEFT_GRAPH[2991], LEFT_GRAPH[2927], LEFT_GRAPH[2863], LEFT_GRAPH[2799], LEFT_GRAPH[2735], LEFT_GRAPH[2671], LEFT_GRAPH[2607]};
					9'd368	:	PATTERN = {LEFT_GRAPH[3056], LEFT_GRAPH[2992], LEFT_GRAPH[2928], LEFT_GRAPH[2864], LEFT_GRAPH[2800], LEFT_GRAPH[2736], LEFT_GRAPH[2672], LEFT_GRAPH[2608]};
					9'd369	:	PATTERN = {LEFT_GRAPH[3057], LEFT_GRAPH[2993], LEFT_GRAPH[2929], LEFT_GRAPH[2865], LEFT_GRAPH[2801], LEFT_GRAPH[2737], LEFT_GRAPH[2673], LEFT_GRAPH[2609]};
					9'd370	:	PATTERN = {LEFT_GRAPH[3058], LEFT_GRAPH[2994], LEFT_GRAPH[2930], LEFT_GRAPH[2866], LEFT_GRAPH[2802], LEFT_GRAPH[2738], LEFT_GRAPH[2674], LEFT_GRAPH[2610]};
					9'd371	:	PATTERN = {LEFT_GRAPH[3059], LEFT_GRAPH[2995], LEFT_GRAPH[2931], LEFT_GRAPH[2867], LEFT_GRAPH[2803], LEFT_GRAPH[2739], LEFT_GRAPH[2675], LEFT_GRAPH[2611]};
					9'd372	:	PATTERN = {LEFT_GRAPH[3060], LEFT_GRAPH[2996], LEFT_GRAPH[2932], LEFT_GRAPH[2868], LEFT_GRAPH[2804], LEFT_GRAPH[2740], LEFT_GRAPH[2676], LEFT_GRAPH[2612]};
					9'd373	:	PATTERN = {LEFT_GRAPH[3061], LEFT_GRAPH[2997], LEFT_GRAPH[2933], LEFT_GRAPH[2869], LEFT_GRAPH[2805], LEFT_GRAPH[2741], LEFT_GRAPH[2677], LEFT_GRAPH[2613]};
					9'd374	:	PATTERN = {LEFT_GRAPH[3062], LEFT_GRAPH[2998], LEFT_GRAPH[2934], LEFT_GRAPH[2870], LEFT_GRAPH[2806], LEFT_GRAPH[2742], LEFT_GRAPH[2678], LEFT_GRAPH[2614]};
					9'd375	:	PATTERN = {LEFT_GRAPH[3063], LEFT_GRAPH[2999], LEFT_GRAPH[2935], LEFT_GRAPH[2871], LEFT_GRAPH[2807], LEFT_GRAPH[2743], LEFT_GRAPH[2679], LEFT_GRAPH[2615]};
					9'd376	:	PATTERN = {LEFT_GRAPH[3064], LEFT_GRAPH[3000], LEFT_GRAPH[2936], LEFT_GRAPH[2872], LEFT_GRAPH[2808], LEFT_GRAPH[2744], LEFT_GRAPH[2680], LEFT_GRAPH[2616]};
					9'd377	:	PATTERN = {LEFT_GRAPH[3065], LEFT_GRAPH[3001], LEFT_GRAPH[2937], LEFT_GRAPH[2873], LEFT_GRAPH[2809], LEFT_GRAPH[2745], LEFT_GRAPH[2681], LEFT_GRAPH[2617]};
					9'd378	:	PATTERN = {LEFT_GRAPH[3066], LEFT_GRAPH[3002], LEFT_GRAPH[2938], LEFT_GRAPH[2874], LEFT_GRAPH[2810], LEFT_GRAPH[2746], LEFT_GRAPH[2682], LEFT_GRAPH[2618]};
					9'd379	:	PATTERN = {LEFT_GRAPH[3067], LEFT_GRAPH[3003], LEFT_GRAPH[2939], LEFT_GRAPH[2875], LEFT_GRAPH[2811], LEFT_GRAPH[2747], LEFT_GRAPH[2683], LEFT_GRAPH[2619]};
					9'd380	:	PATTERN = {LEFT_GRAPH[3068], LEFT_GRAPH[3004], LEFT_GRAPH[2940], LEFT_GRAPH[2876], LEFT_GRAPH[2812], LEFT_GRAPH[2748], LEFT_GRAPH[2684], LEFT_GRAPH[2620]};
					9'd381	:	PATTERN = {LEFT_GRAPH[3069], LEFT_GRAPH[3005], LEFT_GRAPH[2941], LEFT_GRAPH[2877], LEFT_GRAPH[2813], LEFT_GRAPH[2749], LEFT_GRAPH[2685], LEFT_GRAPH[2621]};
					9'd382	:	PATTERN = {LEFT_GRAPH[3070], LEFT_GRAPH[3006], LEFT_GRAPH[2942], LEFT_GRAPH[2878], LEFT_GRAPH[2814], LEFT_GRAPH[2750], LEFT_GRAPH[2686], LEFT_GRAPH[2622]};
					9'd383	:	PATTERN = {LEFT_GRAPH[3071], LEFT_GRAPH[3007], LEFT_GRAPH[2943], LEFT_GRAPH[2879], LEFT_GRAPH[2815], LEFT_GRAPH[2751], LEFT_GRAPH[2687], LEFT_GRAPH[2623]};
					9'd384	:	PATTERN = {LEFT_GRAPH[3520], LEFT_GRAPH[3456], LEFT_GRAPH[3392], LEFT_GRAPH[3328], LEFT_GRAPH[3264], LEFT_GRAPH[3200], LEFT_GRAPH[3136], LEFT_GRAPH[3072]};
					9'd385	:	PATTERN = {LEFT_GRAPH[3521], LEFT_GRAPH[3457], LEFT_GRAPH[3393], LEFT_GRAPH[3329], LEFT_GRAPH[3265], LEFT_GRAPH[3201], LEFT_GRAPH[3137], LEFT_GRAPH[3073]};
					9'd386	:	PATTERN = {LEFT_GRAPH[3522], LEFT_GRAPH[3458], LEFT_GRAPH[3394], LEFT_GRAPH[3330], LEFT_GRAPH[3266], LEFT_GRAPH[3202], LEFT_GRAPH[3138], LEFT_GRAPH[3074]};
					9'd387	:	PATTERN = {LEFT_GRAPH[3523], LEFT_GRAPH[3459], LEFT_GRAPH[3395], LEFT_GRAPH[3331], LEFT_GRAPH[3267], LEFT_GRAPH[3203], LEFT_GRAPH[3139], LEFT_GRAPH[3075]};
					9'd388	:	PATTERN = {LEFT_GRAPH[3524], LEFT_GRAPH[3460], LEFT_GRAPH[3396], LEFT_GRAPH[3332], LEFT_GRAPH[3268], LEFT_GRAPH[3204], LEFT_GRAPH[3140], LEFT_GRAPH[3076]};
					9'd389	:	PATTERN = {LEFT_GRAPH[3525], LEFT_GRAPH[3461], LEFT_GRAPH[3397], LEFT_GRAPH[3333], LEFT_GRAPH[3269], LEFT_GRAPH[3205], LEFT_GRAPH[3141], LEFT_GRAPH[3077]};
					9'd390	:	PATTERN = {LEFT_GRAPH[3526], LEFT_GRAPH[3462], LEFT_GRAPH[3398], LEFT_GRAPH[3334], LEFT_GRAPH[3270], LEFT_GRAPH[3206], LEFT_GRAPH[3142], LEFT_GRAPH[3078]};
					9'd391	:	PATTERN = {LEFT_GRAPH[3527], LEFT_GRAPH[3463], LEFT_GRAPH[3399], LEFT_GRAPH[3335], LEFT_GRAPH[3271], LEFT_GRAPH[3207], LEFT_GRAPH[3143], LEFT_GRAPH[3079]};
					9'd392	:	PATTERN = {LEFT_GRAPH[3528], LEFT_GRAPH[3464], LEFT_GRAPH[3400], LEFT_GRAPH[3336], LEFT_GRAPH[3272], LEFT_GRAPH[3208], LEFT_GRAPH[3144], LEFT_GRAPH[3080]};
					9'd393	:	PATTERN = {LEFT_GRAPH[3529], LEFT_GRAPH[3465], LEFT_GRAPH[3401], LEFT_GRAPH[3337], LEFT_GRAPH[3273], LEFT_GRAPH[3209], LEFT_GRAPH[3145], LEFT_GRAPH[3081]};
					9'd394	:	PATTERN = {LEFT_GRAPH[3530], LEFT_GRAPH[3466], LEFT_GRAPH[3402], LEFT_GRAPH[3338], LEFT_GRAPH[3274], LEFT_GRAPH[3210], LEFT_GRAPH[3146], LEFT_GRAPH[3082]};
					9'd395	:	PATTERN = {LEFT_GRAPH[3531], LEFT_GRAPH[3467], LEFT_GRAPH[3403], LEFT_GRAPH[3339], LEFT_GRAPH[3275], LEFT_GRAPH[3211], LEFT_GRAPH[3147], LEFT_GRAPH[3083]};
					9'd396	:	PATTERN = {LEFT_GRAPH[3532], LEFT_GRAPH[3468], LEFT_GRAPH[3404], LEFT_GRAPH[3340], LEFT_GRAPH[3276], LEFT_GRAPH[3212], LEFT_GRAPH[3148], LEFT_GRAPH[3084]};
					9'd397	:	PATTERN = {LEFT_GRAPH[3533], LEFT_GRAPH[3469], LEFT_GRAPH[3405], LEFT_GRAPH[3341], LEFT_GRAPH[3277], LEFT_GRAPH[3213], LEFT_GRAPH[3149], LEFT_GRAPH[3085]};
					9'd398	:	PATTERN = {LEFT_GRAPH[3534], LEFT_GRAPH[3470], LEFT_GRAPH[3406], LEFT_GRAPH[3342], LEFT_GRAPH[3278], LEFT_GRAPH[3214], LEFT_GRAPH[3150], LEFT_GRAPH[3086]};
					9'd399	:	PATTERN = {LEFT_GRAPH[3535], LEFT_GRAPH[3471], LEFT_GRAPH[3407], LEFT_GRAPH[3343], LEFT_GRAPH[3279], LEFT_GRAPH[3215], LEFT_GRAPH[3151], LEFT_GRAPH[3087]};
					9'd400	:	PATTERN = {LEFT_GRAPH[3536], LEFT_GRAPH[3472], LEFT_GRAPH[3408], LEFT_GRAPH[3344], LEFT_GRAPH[3280], LEFT_GRAPH[3216], LEFT_GRAPH[3152], LEFT_GRAPH[3088]};
					9'd401	:	PATTERN = {LEFT_GRAPH[3537], LEFT_GRAPH[3473], LEFT_GRAPH[3409], LEFT_GRAPH[3345], LEFT_GRAPH[3281], LEFT_GRAPH[3217], LEFT_GRAPH[3153], LEFT_GRAPH[3089]};
					9'd402	:	PATTERN = {LEFT_GRAPH[3538], LEFT_GRAPH[3474], LEFT_GRAPH[3410], LEFT_GRAPH[3346], LEFT_GRAPH[3282], LEFT_GRAPH[3218], LEFT_GRAPH[3154], LEFT_GRAPH[3090]};
					9'd403	:	PATTERN = {LEFT_GRAPH[3539], LEFT_GRAPH[3475], LEFT_GRAPH[3411], LEFT_GRAPH[3347], LEFT_GRAPH[3283], LEFT_GRAPH[3219], LEFT_GRAPH[3155], LEFT_GRAPH[3091]};
					9'd404	:	PATTERN = {LEFT_GRAPH[3540], LEFT_GRAPH[3476], LEFT_GRAPH[3412], LEFT_GRAPH[3348], LEFT_GRAPH[3284], LEFT_GRAPH[3220], LEFT_GRAPH[3156], LEFT_GRAPH[3092]};
					9'd405	:	PATTERN = {LEFT_GRAPH[3541], LEFT_GRAPH[3477], LEFT_GRAPH[3413], LEFT_GRAPH[3349], LEFT_GRAPH[3285], LEFT_GRAPH[3221], LEFT_GRAPH[3157], LEFT_GRAPH[3093]};
					9'd406	:	PATTERN = {LEFT_GRAPH[3542], LEFT_GRAPH[3478], LEFT_GRAPH[3414], LEFT_GRAPH[3350], LEFT_GRAPH[3286], LEFT_GRAPH[3222], LEFT_GRAPH[3158], LEFT_GRAPH[3094]};
					9'd407	:	PATTERN = {LEFT_GRAPH[3543], LEFT_GRAPH[3479], LEFT_GRAPH[3415], LEFT_GRAPH[3351], LEFT_GRAPH[3287], LEFT_GRAPH[3223], LEFT_GRAPH[3159], LEFT_GRAPH[3095]};
					9'd408	:	PATTERN = {LEFT_GRAPH[3544], LEFT_GRAPH[3480], LEFT_GRAPH[3416], LEFT_GRAPH[3352], LEFT_GRAPH[3288], LEFT_GRAPH[3224], LEFT_GRAPH[3160], LEFT_GRAPH[3096]};
					9'd409	:	PATTERN = {LEFT_GRAPH[3545], LEFT_GRAPH[3481], LEFT_GRAPH[3417], LEFT_GRAPH[3353], LEFT_GRAPH[3289], LEFT_GRAPH[3225], LEFT_GRAPH[3161], LEFT_GRAPH[3097]};
					9'd410	:	PATTERN = {LEFT_GRAPH[3546], LEFT_GRAPH[3482], LEFT_GRAPH[3418], LEFT_GRAPH[3354], LEFT_GRAPH[3290], LEFT_GRAPH[3226], LEFT_GRAPH[3162], LEFT_GRAPH[3098]};
					9'd411	:	PATTERN = {LEFT_GRAPH[3547], LEFT_GRAPH[3483], LEFT_GRAPH[3419], LEFT_GRAPH[3355], LEFT_GRAPH[3291], LEFT_GRAPH[3227], LEFT_GRAPH[3163], LEFT_GRAPH[3099]};
					9'd412	:	PATTERN = {LEFT_GRAPH[3548], LEFT_GRAPH[3484], LEFT_GRAPH[3420], LEFT_GRAPH[3356], LEFT_GRAPH[3292], LEFT_GRAPH[3228], LEFT_GRAPH[3164], LEFT_GRAPH[3100]};
					9'd413	:	PATTERN = {LEFT_GRAPH[3549], LEFT_GRAPH[3485], LEFT_GRAPH[3421], LEFT_GRAPH[3357], LEFT_GRAPH[3293], LEFT_GRAPH[3229], LEFT_GRAPH[3165], LEFT_GRAPH[3101]};
					9'd414	:	PATTERN = {LEFT_GRAPH[3550], LEFT_GRAPH[3486], LEFT_GRAPH[3422], LEFT_GRAPH[3358], LEFT_GRAPH[3294], LEFT_GRAPH[3230], LEFT_GRAPH[3166], LEFT_GRAPH[3102]};
					9'd415	:	PATTERN = {LEFT_GRAPH[3551], LEFT_GRAPH[3487], LEFT_GRAPH[3423], LEFT_GRAPH[3359], LEFT_GRAPH[3295], LEFT_GRAPH[3231], LEFT_GRAPH[3167], LEFT_GRAPH[3103]};
					9'd416	:	PATTERN = {LEFT_GRAPH[3552], LEFT_GRAPH[3488], LEFT_GRAPH[3424], LEFT_GRAPH[3360], LEFT_GRAPH[3296], LEFT_GRAPH[3232], LEFT_GRAPH[3168], LEFT_GRAPH[3104]};
					9'd417	:	PATTERN = {LEFT_GRAPH[3553], LEFT_GRAPH[3489], LEFT_GRAPH[3425], LEFT_GRAPH[3361], LEFT_GRAPH[3297], LEFT_GRAPH[3233], LEFT_GRAPH[3169], LEFT_GRAPH[3105]};
					9'd418	:	PATTERN = {LEFT_GRAPH[3554], LEFT_GRAPH[3490], LEFT_GRAPH[3426], LEFT_GRAPH[3362], LEFT_GRAPH[3298], LEFT_GRAPH[3234], LEFT_GRAPH[3170], LEFT_GRAPH[3106]};
					9'd419	:	PATTERN = {LEFT_GRAPH[3555], LEFT_GRAPH[3491], LEFT_GRAPH[3427], LEFT_GRAPH[3363], LEFT_GRAPH[3299], LEFT_GRAPH[3235], LEFT_GRAPH[3171], LEFT_GRAPH[3107]};
					9'd420	:	PATTERN = {LEFT_GRAPH[3556], LEFT_GRAPH[3492], LEFT_GRAPH[3428], LEFT_GRAPH[3364], LEFT_GRAPH[3300], LEFT_GRAPH[3236], LEFT_GRAPH[3172], LEFT_GRAPH[3108]};
					9'd421	:	PATTERN = {LEFT_GRAPH[3557], LEFT_GRAPH[3493], LEFT_GRAPH[3429], LEFT_GRAPH[3365], LEFT_GRAPH[3301], LEFT_GRAPH[3237], LEFT_GRAPH[3173], LEFT_GRAPH[3109]};
					9'd422	:	PATTERN = {LEFT_GRAPH[3558], LEFT_GRAPH[3494], LEFT_GRAPH[3430], LEFT_GRAPH[3366], LEFT_GRAPH[3302], LEFT_GRAPH[3238], LEFT_GRAPH[3174], LEFT_GRAPH[3110]};
					9'd423	:	PATTERN = {LEFT_GRAPH[3559], LEFT_GRAPH[3495], LEFT_GRAPH[3431], LEFT_GRAPH[3367], LEFT_GRAPH[3303], LEFT_GRAPH[3239], LEFT_GRAPH[3175], LEFT_GRAPH[3111]};
					9'd424	:	PATTERN = {LEFT_GRAPH[3560], LEFT_GRAPH[3496], LEFT_GRAPH[3432], LEFT_GRAPH[3368], LEFT_GRAPH[3304], LEFT_GRAPH[3240], LEFT_GRAPH[3176], LEFT_GRAPH[3112]};
					9'd425	:	PATTERN = {LEFT_GRAPH[3561], LEFT_GRAPH[3497], LEFT_GRAPH[3433], LEFT_GRAPH[3369], LEFT_GRAPH[3305], LEFT_GRAPH[3241], LEFT_GRAPH[3177], LEFT_GRAPH[3113]};
					9'd426	:	PATTERN = {LEFT_GRAPH[3562], LEFT_GRAPH[3498], LEFT_GRAPH[3434], LEFT_GRAPH[3370], LEFT_GRAPH[3306], LEFT_GRAPH[3242], LEFT_GRAPH[3178], LEFT_GRAPH[3114]};
					9'd427	:	PATTERN = {LEFT_GRAPH[3563], LEFT_GRAPH[3499], LEFT_GRAPH[3435], LEFT_GRAPH[3371], LEFT_GRAPH[3307], LEFT_GRAPH[3243], LEFT_GRAPH[3179], LEFT_GRAPH[3115]};
					9'd428	:	PATTERN = {LEFT_GRAPH[3564], LEFT_GRAPH[3500], LEFT_GRAPH[3436], LEFT_GRAPH[3372], LEFT_GRAPH[3308], LEFT_GRAPH[3244], LEFT_GRAPH[3180], LEFT_GRAPH[3116]};
					9'd429	:	PATTERN = {LEFT_GRAPH[3565], LEFT_GRAPH[3501], LEFT_GRAPH[3437], LEFT_GRAPH[3373], LEFT_GRAPH[3309], LEFT_GRAPH[3245], LEFT_GRAPH[3181], LEFT_GRAPH[3117]};
					9'd430	:	PATTERN = {LEFT_GRAPH[3566], LEFT_GRAPH[3502], LEFT_GRAPH[3438], LEFT_GRAPH[3374], LEFT_GRAPH[3310], LEFT_GRAPH[3246], LEFT_GRAPH[3182], LEFT_GRAPH[3118]};
					9'd431	:	PATTERN = {LEFT_GRAPH[3567], LEFT_GRAPH[3503], LEFT_GRAPH[3439], LEFT_GRAPH[3375], LEFT_GRAPH[3311], LEFT_GRAPH[3247], LEFT_GRAPH[3183], LEFT_GRAPH[3119]};
					9'd432	:	PATTERN = {LEFT_GRAPH[3568], LEFT_GRAPH[3504], LEFT_GRAPH[3440], LEFT_GRAPH[3376], LEFT_GRAPH[3312], LEFT_GRAPH[3248], LEFT_GRAPH[3184], LEFT_GRAPH[3120]};
					9'd433	:	PATTERN = {LEFT_GRAPH[3569], LEFT_GRAPH[3505], LEFT_GRAPH[3441], LEFT_GRAPH[3377], LEFT_GRAPH[3313], LEFT_GRAPH[3249], LEFT_GRAPH[3185], LEFT_GRAPH[3121]};
					9'd434	:	PATTERN = {LEFT_GRAPH[3570], LEFT_GRAPH[3506], LEFT_GRAPH[3442], LEFT_GRAPH[3378], LEFT_GRAPH[3314], LEFT_GRAPH[3250], LEFT_GRAPH[3186], LEFT_GRAPH[3122]};
					9'd435	:	PATTERN = {LEFT_GRAPH[3571], LEFT_GRAPH[3507], LEFT_GRAPH[3443], LEFT_GRAPH[3379], LEFT_GRAPH[3315], LEFT_GRAPH[3251], LEFT_GRAPH[3187], LEFT_GRAPH[3123]};
					9'd436	:	PATTERN = {LEFT_GRAPH[3572], LEFT_GRAPH[3508], LEFT_GRAPH[3444], LEFT_GRAPH[3380], LEFT_GRAPH[3316], LEFT_GRAPH[3252], LEFT_GRAPH[3188], LEFT_GRAPH[3124]};
					9'd437	:	PATTERN = {LEFT_GRAPH[3573], LEFT_GRAPH[3509], LEFT_GRAPH[3445], LEFT_GRAPH[3381], LEFT_GRAPH[3317], LEFT_GRAPH[3253], LEFT_GRAPH[3189], LEFT_GRAPH[3125]};
					9'd438	:	PATTERN = {LEFT_GRAPH[3574], LEFT_GRAPH[3510], LEFT_GRAPH[3446], LEFT_GRAPH[3382], LEFT_GRAPH[3318], LEFT_GRAPH[3254], LEFT_GRAPH[3190], LEFT_GRAPH[3126]};
					9'd439	:	PATTERN = {LEFT_GRAPH[3575], LEFT_GRAPH[3511], LEFT_GRAPH[3447], LEFT_GRAPH[3383], LEFT_GRAPH[3319], LEFT_GRAPH[3255], LEFT_GRAPH[3191], LEFT_GRAPH[3127]};
					9'd440	:	PATTERN = {LEFT_GRAPH[3576], LEFT_GRAPH[3512], LEFT_GRAPH[3448], LEFT_GRAPH[3384], LEFT_GRAPH[3320], LEFT_GRAPH[3256], LEFT_GRAPH[3192], LEFT_GRAPH[3128]};
					9'd441	:	PATTERN = {LEFT_GRAPH[3577], LEFT_GRAPH[3513], LEFT_GRAPH[3449], LEFT_GRAPH[3385], LEFT_GRAPH[3321], LEFT_GRAPH[3257], LEFT_GRAPH[3193], LEFT_GRAPH[3129]};
					9'd442	:	PATTERN = {LEFT_GRAPH[3578], LEFT_GRAPH[3514], LEFT_GRAPH[3450], LEFT_GRAPH[3386], LEFT_GRAPH[3322], LEFT_GRAPH[3258], LEFT_GRAPH[3194], LEFT_GRAPH[3130]};
					9'd443	:	PATTERN = {LEFT_GRAPH[3579], LEFT_GRAPH[3515], LEFT_GRAPH[3451], LEFT_GRAPH[3387], LEFT_GRAPH[3323], LEFT_GRAPH[3259], LEFT_GRAPH[3195], LEFT_GRAPH[3131]};
					9'd444	:	PATTERN = {LEFT_GRAPH[3580], LEFT_GRAPH[3516], LEFT_GRAPH[3452], LEFT_GRAPH[3388], LEFT_GRAPH[3324], LEFT_GRAPH[3260], LEFT_GRAPH[3196], LEFT_GRAPH[3132]};
					9'd445	:	PATTERN = {LEFT_GRAPH[3581], LEFT_GRAPH[3517], LEFT_GRAPH[3453], LEFT_GRAPH[3389], LEFT_GRAPH[3325], LEFT_GRAPH[3261], LEFT_GRAPH[3197], LEFT_GRAPH[3133]};
					9'd446	:	PATTERN = {LEFT_GRAPH[3582], LEFT_GRAPH[3518], LEFT_GRAPH[3454], LEFT_GRAPH[3390], LEFT_GRAPH[3326], LEFT_GRAPH[3262], LEFT_GRAPH[3198], LEFT_GRAPH[3134]};
					9'd447	:	PATTERN = {LEFT_GRAPH[3583], LEFT_GRAPH[3519], LEFT_GRAPH[3455], LEFT_GRAPH[3391], LEFT_GRAPH[3327], LEFT_GRAPH[3263], LEFT_GRAPH[3199], LEFT_GRAPH[3135]};
					9'd448	:	PATTERN = {LEFT_GRAPH[4032], LEFT_GRAPH[3968], LEFT_GRAPH[3904], LEFT_GRAPH[3840], LEFT_GRAPH[3776], LEFT_GRAPH[3712], LEFT_GRAPH[3648], LEFT_GRAPH[3584]};
					9'd449	:	PATTERN = {LEFT_GRAPH[4033], LEFT_GRAPH[3969], LEFT_GRAPH[3905], LEFT_GRAPH[3841], LEFT_GRAPH[3777], LEFT_GRAPH[3713], LEFT_GRAPH[3649], LEFT_GRAPH[3585]};
					9'd450	:	PATTERN = {LEFT_GRAPH[4034], LEFT_GRAPH[3970], LEFT_GRAPH[3906], LEFT_GRAPH[3842], LEFT_GRAPH[3778], LEFT_GRAPH[3714], LEFT_GRAPH[3650], LEFT_GRAPH[3586]};
					9'd451	:	PATTERN = {LEFT_GRAPH[4035], LEFT_GRAPH[3971], LEFT_GRAPH[3907], LEFT_GRAPH[3843], LEFT_GRAPH[3779], LEFT_GRAPH[3715], LEFT_GRAPH[3651], LEFT_GRAPH[3587]};
					9'd452	:	PATTERN = {LEFT_GRAPH[4036], LEFT_GRAPH[3972], LEFT_GRAPH[3908], LEFT_GRAPH[3844], LEFT_GRAPH[3780], LEFT_GRAPH[3716], LEFT_GRAPH[3652], LEFT_GRAPH[3588]};
					9'd453	:	PATTERN = {LEFT_GRAPH[4037], LEFT_GRAPH[3973], LEFT_GRAPH[3909], LEFT_GRAPH[3845], LEFT_GRAPH[3781], LEFT_GRAPH[3717], LEFT_GRAPH[3653], LEFT_GRAPH[3589]};
					9'd454	:	PATTERN = {LEFT_GRAPH[4038], LEFT_GRAPH[3974], LEFT_GRAPH[3910], LEFT_GRAPH[3846], LEFT_GRAPH[3782], LEFT_GRAPH[3718], LEFT_GRAPH[3654], LEFT_GRAPH[3590]};
					9'd455	:	PATTERN = {LEFT_GRAPH[4039], LEFT_GRAPH[3975], LEFT_GRAPH[3911], LEFT_GRAPH[3847], LEFT_GRAPH[3783], LEFT_GRAPH[3719], LEFT_GRAPH[3655], LEFT_GRAPH[3591]};
					9'd456	:	PATTERN = {LEFT_GRAPH[4040], LEFT_GRAPH[3976], LEFT_GRAPH[3912], LEFT_GRAPH[3848], LEFT_GRAPH[3784], LEFT_GRAPH[3720], LEFT_GRAPH[3656], LEFT_GRAPH[3592]};
					9'd457	:	PATTERN = {LEFT_GRAPH[4041], LEFT_GRAPH[3977], LEFT_GRAPH[3913], LEFT_GRAPH[3849], LEFT_GRAPH[3785], LEFT_GRAPH[3721], LEFT_GRAPH[3657], LEFT_GRAPH[3593]};
					9'd458	:	PATTERN = {LEFT_GRAPH[4042], LEFT_GRAPH[3978], LEFT_GRAPH[3914], LEFT_GRAPH[3850], LEFT_GRAPH[3786], LEFT_GRAPH[3722], LEFT_GRAPH[3658], LEFT_GRAPH[3594]};
					9'd459	:	PATTERN = {LEFT_GRAPH[4043], LEFT_GRAPH[3979], LEFT_GRAPH[3915], LEFT_GRAPH[3851], LEFT_GRAPH[3787], LEFT_GRAPH[3723], LEFT_GRAPH[3659], LEFT_GRAPH[3595]};
					9'd460	:	PATTERN = {LEFT_GRAPH[4044], LEFT_GRAPH[3980], LEFT_GRAPH[3916], LEFT_GRAPH[3852], LEFT_GRAPH[3788], LEFT_GRAPH[3724], LEFT_GRAPH[3660], LEFT_GRAPH[3596]};
					9'd461	:	PATTERN = {LEFT_GRAPH[4045], LEFT_GRAPH[3981], LEFT_GRAPH[3917], LEFT_GRAPH[3853], LEFT_GRAPH[3789], LEFT_GRAPH[3725], LEFT_GRAPH[3661], LEFT_GRAPH[3597]};
					9'd462	:	PATTERN = {LEFT_GRAPH[4046], LEFT_GRAPH[3982], LEFT_GRAPH[3918], LEFT_GRAPH[3854], LEFT_GRAPH[3790], LEFT_GRAPH[3726], LEFT_GRAPH[3662], LEFT_GRAPH[3598]};
					9'd463	:	PATTERN = {LEFT_GRAPH[4047], LEFT_GRAPH[3983], LEFT_GRAPH[3919], LEFT_GRAPH[3855], LEFT_GRAPH[3791], LEFT_GRAPH[3727], LEFT_GRAPH[3663], LEFT_GRAPH[3599]};
					9'd464	:	PATTERN = {LEFT_GRAPH[4048], LEFT_GRAPH[3984], LEFT_GRAPH[3920], LEFT_GRAPH[3856], LEFT_GRAPH[3792], LEFT_GRAPH[3728], LEFT_GRAPH[3664], LEFT_GRAPH[3600]};
					9'd465	:	PATTERN = {LEFT_GRAPH[4049], LEFT_GRAPH[3985], LEFT_GRAPH[3921], LEFT_GRAPH[3857], LEFT_GRAPH[3793], LEFT_GRAPH[3729], LEFT_GRAPH[3665], LEFT_GRAPH[3601]};
					9'd466	:	PATTERN = {LEFT_GRAPH[4050], LEFT_GRAPH[3986], LEFT_GRAPH[3922], LEFT_GRAPH[3858], LEFT_GRAPH[3794], LEFT_GRAPH[3730], LEFT_GRAPH[3666], LEFT_GRAPH[3602]};
					9'd467	:	PATTERN = {LEFT_GRAPH[4051], LEFT_GRAPH[3987], LEFT_GRAPH[3923], LEFT_GRAPH[3859], LEFT_GRAPH[3795], LEFT_GRAPH[3731], LEFT_GRAPH[3667], LEFT_GRAPH[3603]};
					9'd468	:	PATTERN = {LEFT_GRAPH[4052], LEFT_GRAPH[3988], LEFT_GRAPH[3924], LEFT_GRAPH[3860], LEFT_GRAPH[3796], LEFT_GRAPH[3732], LEFT_GRAPH[3668], LEFT_GRAPH[3604]};
					9'd469	:	PATTERN = {LEFT_GRAPH[4053], LEFT_GRAPH[3989], LEFT_GRAPH[3925], LEFT_GRAPH[3861], LEFT_GRAPH[3797], LEFT_GRAPH[3733], LEFT_GRAPH[3669], LEFT_GRAPH[3605]};
					9'd470	:	PATTERN = {LEFT_GRAPH[4054], LEFT_GRAPH[3990], LEFT_GRAPH[3926], LEFT_GRAPH[3862], LEFT_GRAPH[3798], LEFT_GRAPH[3734], LEFT_GRAPH[3670], LEFT_GRAPH[3606]};
					9'd471	:	PATTERN = {LEFT_GRAPH[4055], LEFT_GRAPH[3991], LEFT_GRAPH[3927], LEFT_GRAPH[3863], LEFT_GRAPH[3799], LEFT_GRAPH[3735], LEFT_GRAPH[3671], LEFT_GRAPH[3607]};
					9'd472	:	PATTERN = {LEFT_GRAPH[4056], LEFT_GRAPH[3992], LEFT_GRAPH[3928], LEFT_GRAPH[3864], LEFT_GRAPH[3800], LEFT_GRAPH[3736], LEFT_GRAPH[3672], LEFT_GRAPH[3608]};
					9'd473	:	PATTERN = {LEFT_GRAPH[4057], LEFT_GRAPH[3993], LEFT_GRAPH[3929], LEFT_GRAPH[3865], LEFT_GRAPH[3801], LEFT_GRAPH[3737], LEFT_GRAPH[3673], LEFT_GRAPH[3609]};
					9'd474	:	PATTERN = {LEFT_GRAPH[4058], LEFT_GRAPH[3994], LEFT_GRAPH[3930], LEFT_GRAPH[3866], LEFT_GRAPH[3802], LEFT_GRAPH[3738], LEFT_GRAPH[3674], LEFT_GRAPH[3610]};
					9'd475	:	PATTERN = {LEFT_GRAPH[4059], LEFT_GRAPH[3995], LEFT_GRAPH[3931], LEFT_GRAPH[3867], LEFT_GRAPH[3803], LEFT_GRAPH[3739], LEFT_GRAPH[3675], LEFT_GRAPH[3611]};
					9'd476	:	PATTERN = {LEFT_GRAPH[4060], LEFT_GRAPH[3996], LEFT_GRAPH[3932], LEFT_GRAPH[3868], LEFT_GRAPH[3804], LEFT_GRAPH[3740], LEFT_GRAPH[3676], LEFT_GRAPH[3612]};
					9'd477	:	PATTERN = {LEFT_GRAPH[4061], LEFT_GRAPH[3997], LEFT_GRAPH[3933], LEFT_GRAPH[3869], LEFT_GRAPH[3805], LEFT_GRAPH[3741], LEFT_GRAPH[3677], LEFT_GRAPH[3613]};
					9'd478	:	PATTERN = {LEFT_GRAPH[4062], LEFT_GRAPH[3998], LEFT_GRAPH[3934], LEFT_GRAPH[3870], LEFT_GRAPH[3806], LEFT_GRAPH[3742], LEFT_GRAPH[3678], LEFT_GRAPH[3614]};
					9'd479	:	PATTERN = {LEFT_GRAPH[4063], LEFT_GRAPH[3999], LEFT_GRAPH[3935], LEFT_GRAPH[3871], LEFT_GRAPH[3807], LEFT_GRAPH[3743], LEFT_GRAPH[3679], LEFT_GRAPH[3615]};
					9'd480	:	PATTERN = {LEFT_GRAPH[4064], LEFT_GRAPH[4000], LEFT_GRAPH[3936], LEFT_GRAPH[3872], LEFT_GRAPH[3808], LEFT_GRAPH[3744], LEFT_GRAPH[3680], LEFT_GRAPH[3616]};
					9'd481	:	PATTERN = {LEFT_GRAPH[4065], LEFT_GRAPH[4001], LEFT_GRAPH[3937], LEFT_GRAPH[3873], LEFT_GRAPH[3809], LEFT_GRAPH[3745], LEFT_GRAPH[3681], LEFT_GRAPH[3617]};
					9'd482	:	PATTERN = {LEFT_GRAPH[4066], LEFT_GRAPH[4002], LEFT_GRAPH[3938], LEFT_GRAPH[3874], LEFT_GRAPH[3810], LEFT_GRAPH[3746], LEFT_GRAPH[3682], LEFT_GRAPH[3618]};
					9'd483	:	PATTERN = {LEFT_GRAPH[4067], LEFT_GRAPH[4003], LEFT_GRAPH[3939], LEFT_GRAPH[3875], LEFT_GRAPH[3811], LEFT_GRAPH[3747], LEFT_GRAPH[3683], LEFT_GRAPH[3619]};
					9'd484	:	PATTERN = {LEFT_GRAPH[4068], LEFT_GRAPH[4004], LEFT_GRAPH[3940], LEFT_GRAPH[3876], LEFT_GRAPH[3812], LEFT_GRAPH[3748], LEFT_GRAPH[3684], LEFT_GRAPH[3620]};
					9'd485	:	PATTERN = {LEFT_GRAPH[4069], LEFT_GRAPH[4005], LEFT_GRAPH[3941], LEFT_GRAPH[3877], LEFT_GRAPH[3813], LEFT_GRAPH[3749], LEFT_GRAPH[3685], LEFT_GRAPH[3621]};
					9'd486	:	PATTERN = {LEFT_GRAPH[4070], LEFT_GRAPH[4006], LEFT_GRAPH[3942], LEFT_GRAPH[3878], LEFT_GRAPH[3814], LEFT_GRAPH[3750], LEFT_GRAPH[3686], LEFT_GRAPH[3622]};
					9'd487	:	PATTERN = {LEFT_GRAPH[4071], LEFT_GRAPH[4007], LEFT_GRAPH[3943], LEFT_GRAPH[3879], LEFT_GRAPH[3815], LEFT_GRAPH[3751], LEFT_GRAPH[3687], LEFT_GRAPH[3623]};
					9'd488	:	PATTERN = {LEFT_GRAPH[4072], LEFT_GRAPH[4008], LEFT_GRAPH[3944], LEFT_GRAPH[3880], LEFT_GRAPH[3816], LEFT_GRAPH[3752], LEFT_GRAPH[3688], LEFT_GRAPH[3624]};
					9'd489	:	PATTERN = {LEFT_GRAPH[4073], LEFT_GRAPH[4009], LEFT_GRAPH[3945], LEFT_GRAPH[3881], LEFT_GRAPH[3817], LEFT_GRAPH[3753], LEFT_GRAPH[3689], LEFT_GRAPH[3625]};
					9'd490	:	PATTERN = {LEFT_GRAPH[4074], LEFT_GRAPH[4010], LEFT_GRAPH[3946], LEFT_GRAPH[3882], LEFT_GRAPH[3818], LEFT_GRAPH[3754], LEFT_GRAPH[3690], LEFT_GRAPH[3626]};
					9'd491	:	PATTERN = {LEFT_GRAPH[4075], LEFT_GRAPH[4011], LEFT_GRAPH[3947], LEFT_GRAPH[3883], LEFT_GRAPH[3819], LEFT_GRAPH[3755], LEFT_GRAPH[3691], LEFT_GRAPH[3627]};
					9'd492	:	PATTERN = {LEFT_GRAPH[4076], LEFT_GRAPH[4012], LEFT_GRAPH[3948], LEFT_GRAPH[3884], LEFT_GRAPH[3820], LEFT_GRAPH[3756], LEFT_GRAPH[3692], LEFT_GRAPH[3628]};
					9'd493	:	PATTERN = {LEFT_GRAPH[4077], LEFT_GRAPH[4013], LEFT_GRAPH[3949], LEFT_GRAPH[3885], LEFT_GRAPH[3821], LEFT_GRAPH[3757], LEFT_GRAPH[3693], LEFT_GRAPH[3629]};
					9'd494	:	PATTERN = {LEFT_GRAPH[4078], LEFT_GRAPH[4014], LEFT_GRAPH[3950], LEFT_GRAPH[3886], LEFT_GRAPH[3822], LEFT_GRAPH[3758], LEFT_GRAPH[3694], LEFT_GRAPH[3630]};
					9'd495	:	PATTERN = {LEFT_GRAPH[4079], LEFT_GRAPH[4015], LEFT_GRAPH[3951], LEFT_GRAPH[3887], LEFT_GRAPH[3823], LEFT_GRAPH[3759], LEFT_GRAPH[3695], LEFT_GRAPH[3631]};
					9'd496	:	PATTERN = {LEFT_GRAPH[4080], LEFT_GRAPH[4016], LEFT_GRAPH[3952], LEFT_GRAPH[3888], LEFT_GRAPH[3824], LEFT_GRAPH[3760], LEFT_GRAPH[3696], LEFT_GRAPH[3632]};
					9'd497	:	PATTERN = {LEFT_GRAPH[4081], LEFT_GRAPH[4017], LEFT_GRAPH[3953], LEFT_GRAPH[3889], LEFT_GRAPH[3825], LEFT_GRAPH[3761], LEFT_GRAPH[3697], LEFT_GRAPH[3633]};
					9'd498	:	PATTERN = {LEFT_GRAPH[4082], LEFT_GRAPH[4018], LEFT_GRAPH[3954], LEFT_GRAPH[3890], LEFT_GRAPH[3826], LEFT_GRAPH[3762], LEFT_GRAPH[3698], LEFT_GRAPH[3634]};
					9'd499	:	PATTERN = {LEFT_GRAPH[4083], LEFT_GRAPH[4019], LEFT_GRAPH[3955], LEFT_GRAPH[3891], LEFT_GRAPH[3827], LEFT_GRAPH[3763], LEFT_GRAPH[3699], LEFT_GRAPH[3635]};
					9'd500	:	PATTERN = {LEFT_GRAPH[4084], LEFT_GRAPH[4020], LEFT_GRAPH[3956], LEFT_GRAPH[3892], LEFT_GRAPH[3828], LEFT_GRAPH[3764], LEFT_GRAPH[3700], LEFT_GRAPH[3636]};
					9'd501	:	PATTERN = {LEFT_GRAPH[4085], LEFT_GRAPH[4021], LEFT_GRAPH[3957], LEFT_GRAPH[3893], LEFT_GRAPH[3829], LEFT_GRAPH[3765], LEFT_GRAPH[3701], LEFT_GRAPH[3637]};
					9'd502	:	PATTERN = {LEFT_GRAPH[4086], LEFT_GRAPH[4022], LEFT_GRAPH[3958], LEFT_GRAPH[3894], LEFT_GRAPH[3830], LEFT_GRAPH[3766], LEFT_GRAPH[3702], LEFT_GRAPH[3638]};
					9'd503	:	PATTERN = {LEFT_GRAPH[4087], LEFT_GRAPH[4023], LEFT_GRAPH[3959], LEFT_GRAPH[3895], LEFT_GRAPH[3831], LEFT_GRAPH[3767], LEFT_GRAPH[3703], LEFT_GRAPH[3639]};
					9'd504	:	PATTERN = {LEFT_GRAPH[4088], LEFT_GRAPH[4024], LEFT_GRAPH[3960], LEFT_GRAPH[3896], LEFT_GRAPH[3832], LEFT_GRAPH[3768], LEFT_GRAPH[3704], LEFT_GRAPH[3640]};
					9'd505	:	PATTERN = {LEFT_GRAPH[4089], LEFT_GRAPH[4025], LEFT_GRAPH[3961], LEFT_GRAPH[3897], LEFT_GRAPH[3833], LEFT_GRAPH[3769], LEFT_GRAPH[3705], LEFT_GRAPH[3641]};
					9'd506	:	PATTERN = {LEFT_GRAPH[4090], LEFT_GRAPH[4026], LEFT_GRAPH[3962], LEFT_GRAPH[3898], LEFT_GRAPH[3834], LEFT_GRAPH[3770], LEFT_GRAPH[3706], LEFT_GRAPH[3642]};
					9'd507	:	PATTERN = {LEFT_GRAPH[4091], LEFT_GRAPH[4027], LEFT_GRAPH[3963], LEFT_GRAPH[3899], LEFT_GRAPH[3835], LEFT_GRAPH[3771], LEFT_GRAPH[3707], LEFT_GRAPH[3643]};
					9'd508	:	PATTERN = {LEFT_GRAPH[4092], LEFT_GRAPH[4028], LEFT_GRAPH[3964], LEFT_GRAPH[3900], LEFT_GRAPH[3836], LEFT_GRAPH[3772], LEFT_GRAPH[3708], LEFT_GRAPH[3644]};
					9'd509	:	PATTERN = {LEFT_GRAPH[4093], LEFT_GRAPH[4029], LEFT_GRAPH[3965], LEFT_GRAPH[3901], LEFT_GRAPH[3837], LEFT_GRAPH[3773], LEFT_GRAPH[3709], LEFT_GRAPH[3645]};
					9'd510	:	PATTERN = {LEFT_GRAPH[4094], LEFT_GRAPH[4030], LEFT_GRAPH[3966], LEFT_GRAPH[3902], LEFT_GRAPH[3838], LEFT_GRAPH[3774], LEFT_GRAPH[3710], LEFT_GRAPH[3646]};
					9'd511	:	PATTERN = {LEFT_GRAPH[4095], LEFT_GRAPH[4031], LEFT_GRAPH[3967], LEFT_GRAPH[3903], LEFT_GRAPH[3839], LEFT_GRAPH[3775], LEFT_GRAPH[3711], LEFT_GRAPH[3647]};
				endcase
			endcase
	endcase
  end

endmodule
