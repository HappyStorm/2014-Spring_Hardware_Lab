`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:32:26 06/23/2014 
// Design Name: 
// Module Name:    TAIKO_CONTROL 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module TAIKO_CONTROL(GL, GR, score_tens, score_unit, Melody, pre_Melody, pp_Melody, ppp_Melody, pppp_Melody, KEY_IN, press, isfinish, valid, reset, clk_1Hz, clk_10Hz, clk_100Hz, clk_500ms, clk_100KHz, clk_1s ,clk_1us, clk);
	
	input reset, clk_1Hz, clk_10Hz, clk_100Hz, clk_500ms, clk_100KHz, clk_1s, clk_1us, clk;
	input valid;
	input [4:0] Melody;
	input [4:0] pre_Melody;
	input [4:0] pp_Melody;
	input [4:0] ppp_Melody;
	input [4:0] pppp_Melody;
	input [4:0] KEY_IN;
	input press;
	input isfinish;
	
	output reg [3:0] score_tens;
	output reg [3:0] score_unit;
	output reg [0:4095] GL;
	output reg [0:4095] GR;
	
	reg [1:0] state;
	reg [3:0] tmp_score_tens = 4'b 0;
	reg [3:0] tmp_score_unit = 4'b 0;
	reg  flag_state = 0;
	reg  flag_point = 0;
	
//	reg [4:0] tmp_melody = 0;
//	wire [4:0] tmp_melody;
	
	// Check if the input equals to the melody, if yes, score++, if not, do nothing
//	always @(posedge clk_1s or negedge reset) begin
//		if(!reset) begin
//			tmp_score_tens <= 0;
//			tmp_score_unit <= 0;
//		end
//		else begin 
//			if(valid) begin
//				if(KEY_IN==Melody) begin
//					if(tmp_score_unit==9) begin
//						tmp_score_tens <= (tmp_score_tens+1);
//						tmp_score_unit <= 0;
//					end
//					else begin
//						tmp_score_unit <= (tmp_score_unit+1);
//					end
//				end
//				else begin
//				end
//			end
//			else begin
//			end
//		end
//	end
	
	
	always @(posedge clk_1s or negedge reset) begin	// 0: �S��	1:����	(state = 1: hit)	(state = 2: miss)
//		tmp_melody = Melody;
		if(!press || !reset) begin
			if(!reset) begin
				score_tens <= 0;
				score_unit <= 0;
			end
			else begin
			end
			state <= 2'b00;
			flag_state <= 0;
		end
		else begin
			score_tens <= tmp_score_tens;
			score_unit <= tmp_score_unit;
			if(KEY_IN==pppp_Melody) begin
				if(flag_state==0) begin
					state <= 2'b01;
					flag_state <= 1;
				end
				else begin
				end
			end
			else begin
				if(flag_state==0) begin
					state <= 2'b10;
					flag_state <= 1;
				end
				else begin
				end
			end
		end
	end
//	assign tmp_melody = Melody;
	
	always @(posedge clk_1s) begin
		if(valid) begin	
			if(KEY_IN==pppp_Melody) begin
				if(flag_point==0) begin
					if(score_unit==9) begin
						tmp_score_tens <= (score_tens+1);
						tmp_score_unit <= 0;
					end
					else begin
						tmp_score_tens <= score_tens;
						tmp_score_unit <= (score_unit+1);
					end
					flag_point <= 1;
				end
				else begin
				end
				
				
			end
			else begin
				flag_point <= 0;
			end
		end
		else begin
			tmp_score_tens <= 4'b 0;
			tmp_score_unit <= 4'b 0;
		end
	end
	
//	always @(posedge clk_1s or negedge reset) begin	// 0: �S��	1:����	(state = 1: hit)	(state = 2: miss)
//		if(!press || !reset) begin
//			state <= 2'b00;
//				GR[   0:  63] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[  64: 127] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 128: 191] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 192: 255] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 256: 319] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 320: 383] <= 64'b1011101110111011101110111011101110111011101110111011101110111011;
//				GR[ 384: 447] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
//				GR[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 704: 767] <= 64'b0000111111100111111100111111000000000000000000000000000000000000;
//				GR[ 768: 831] <= 64'b0000000100000100000100100001000000000000000000000000000000000000;
//				GR[ 832: 895] <= 64'b0000000100000100000100100001000000000000000000000000000000000000;
//				GR[ 896: 959] <= 64'b0000000100000100000100100001000000000000000000000000000000000000;
//				GR[ 960:1023] <= 64'b0000000100000111111100111111000000000000000000000000000000000000;
//				GR[1024:1087] <= 64'b0000000100000100000100100000000000000000000000000000000000000000;
//				GR[1088:1151] <= 64'b0000000100000100000100100000000000000000000000000000000000000000;
//				GR[1152:1215] <= 64'b0000000100000100000100100000000000000000000000000000000000000000;
//				GR[1216:1279] <= 64'b0000000100000100000100100000000000000000000000000000000000000000;
//				GR[1280:1343] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1344:1407] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1408:1471] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1472:1535] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1536:1599] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1600:1663] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1664:1727] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1728:1791] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1792:1855] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1856:1919] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1920:1983] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1984:2047] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[2048:2111] <= 64'b0000000000000000000000000000000000111111000000011000000000000000;
//				GR[2112:2175] <= 64'b0000000000000000000000000000000000111111000000011000000000000000;
//				GR[2176:2239] <= 64'b0000000000000000000000000000000000000000000000011000000000000000;
//				GR[2240:2303] <= 64'b0000000000000000000000000000000000000000000000011000000000000000;
//				GR[2304:2367] <= 64'b0000000000000000000000000000000000001100000011111111100000000000;
//				GR[2368:2431] <= 64'b0000000000000000000000000000000000001100000011111111100000000000;
//				GR[2432:2495] <= 64'b0000000000000000000000000000000000001100000000011000000000000000;
//				GR[2496:2559] <= 64'b0000000000000000000000000000000000001100000000011000000000000000;
//				GR[2560:2623] <= 64'b0000000000000000000000000000000000001100000000011000000000000000;
//				GR[2624:2687] <= 64'b0000000000000000000000000000000000001100000000011000000000000000;
//				GR[2688:2751] <= 64'b0000000000000000000000000000000000001100000000011001100000000000;
//				GR[2752:2815] <= 64'b0000000000000000000000000000000000001100000000011001100000000000;
//				GR[2816:2879] <= 64'b0000000000000000000000000000000000001100000000011111100000000000;
//				GR[2880:2943] <= 64'b0000000000000000000000000000000000001100000000011111100000000000;
//				GR[2944:3007] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3008:3071] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3072:3135] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3136:3199] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3584:3647] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
//				GR[3648:3711] <= 64'b1110111011101110111011101110111011101110111011101110111011101110;
//				GR[3712:3775] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3776:3839] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3840:3903] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3904:3967] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3968:4031] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[4032:4095] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//		end
//		else begin
//			if(KEY_IN==Melody) begin
//				state <= 2'b01;
//				GR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[  64: 127] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 128: 191] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 192: 255] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 256: 319] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
//				GR[ 320: 383] <= 64'b1010101010101010101010101010101010101010101010101010101010101010;
//				GR[ 384: 447] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
//				GR[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 832: 895] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 896: 959] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 960:1023] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1024:1087] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[1088:1151] <= 64'b0000000001000000000000010000000111111000000111111111111111000000;
//				GR[1152:1215] <= 64'b0000000001000000000000010000000111111000000000000010000000000000;
//				GR[1216:1279] <= 64'b0000000001000000000000010000000111111000000000000010000000000000;
//				GR[1280:1343] <= 64'b0000000001000000000000010000000111111000000000000010000000000000;
//				GR[1344:1407] <= 64'b0000000001000000000000010000000111111000000000000010000000000000;
//				GR[1408:1471] <= 64'b0000000001000000000000010000000111111000000000000010000000000000;
//				GR[1472:1535] <= 64'b0000000001000000000000010000000000000000000000000010000000000000;
//				GR[1536:1599] <= 64'b0000000001000000000000010000000000000000000000000010000000000000;
//				GR[1600:1663] <= 64'b0000000001000000000000010000000000000000000000000010000000000000;
//				GR[1664:1727] <= 64'b0000000001000000000000010000000000000000000000000010000000000000;
//				GR[1728:1791] <= 64'b0000000001000000000000010000000000000000000000000010000000000000;
//				GR[1792:1855] <= 64'b0000000001000000000000010000000000000000000000000010000000000000;
//				GR[1856:1919] <= 64'b0000000001000000000000010000000000000000000000000010000000000000;
//				GR[1920:1983] <= 64'b0000000001111111111111110000000111111000000000000010000000000000;
//				GR[1984:2047] <= 64'b0000000001000000000000010000000110001000000000000010000000000000;
//				GR[2048:2111] <= 64'b0000000001000000000000010000000101001000000000000010000000000000;
//				GR[2112:2175] <= 64'b0000000001000000000000010000000100101000000000000010000000000000;
//				GR[2176:2239] <= 64'b0000000001000000000000010000000100011000000000000010000000000000;
//				GR[2240:2303] <= 64'b0000000001000000000000010000000100101000000000000010000000000000;
//				GR[2304:2367] <= 64'b0000000001000000000000010000000101001000000000000010000000000000;
//				GR[2368:2431] <= 64'b0000000001000000000000010000000110001000000000000010000000000000;
//				GR[2432:2495] <= 64'b0000000001000000000000010000000101001000000000000010000000000000;
//				GR[2496:2559] <= 64'b0000000001000000000000010000000100101000000000000010000000000000;
//				GR[2560:2623] <= 64'b0000000001000000000000010000000100011000000000000010000000000000;
//				GR[2624:2687] <= 64'b0000000001000000000000010000000100101000000000000010000000000000;
//				GR[2688:2751] <= 64'b0000000001000000000000010000000101001000000000000010000000000000;
//				GR[2752:2815] <= 64'b0000000001000000000000010000000110001000000000000010000000000000;
//				GR[2816:2879] <= 64'b0000000001000000000000010000000111111000000000000010000000000000;
//				GR[2880:2943] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[2944:3007] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3008:3071] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3072:3135] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3136:3199] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3584:3647] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
//				GR[3648:3711] <= 64'b1010101010101010101010101010101010101010101010101010101010101010;
//				GR[3712:3775] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
//				GR[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//			end
//			else begin
//				state <= 2'b10;
//				GR[   0:  63] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[  64: 127] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 128: 191] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 192: 255] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 256: 319] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[ 320: 383] <= 64'b1011101110111011101110111011101110111011101110111011101110111011;
//				GR[ 384: 447] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
//				GR[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 832: 895] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[ 896: 959] <= 64'b0001000000000000000000000111111111000001111111110000111111111000;
//				GR[ 960:1023] <= 64'b0001000000000000000000000111111111000001000000010000100000001000;
//				GR[1024:1087] <= 64'b0001000000000000000000000111111111000001000000010000100000001000;
//				GR[1088:1151] <= 64'b0001111111111111110000000111111111000001000000010000100000001000;
//				GR[1152:1215] <= 64'b0001000000100000010000000111111111000001000000010000100000001000;
//				GR[1216:1279] <= 64'b0001000000100000010000000111111111000001000000000000100000000000;
//				GR[1280:1343] <= 64'b0001000000100000010000000111111111000001000000000000100000000000;
//				GR[1344:1407] <= 64'b0001000000100000010000000000000000000001000000000000100000000000;
//				GR[1408:1471] <= 64'b0001000000100000010000000000000000000001000000000000100000000000;
//				GR[1472:1535] <= 64'b0001000000100000010000000000000000000001000000000000100000000000;
//				GR[1536:1599] <= 64'b0001000000100000010000000000000000000001000000000000100000000000;
//				GR[1600:1663] <= 64'b0001000000100000010000000111111111000001000000000000100000000000;
//				GR[1664:1727] <= 64'b0001000000100000010000000100000011000001000000000000100000000000;
//				GR[1728:1791] <= 64'b0001000000100000010000000100000101000001000000000000100000000000;
//				GR[1792:1855] <= 64'b0001000000100000010000000100001001000001000000000000100000000000;
//				GR[1856:1919] <= 64'b0001000000100000010000000100010001000001111111110000111111111000;
//				GR[1920:1983] <= 64'b0001000000100000010000000100100001000000000000010000000000001000;
//				GR[1984:2047] <= 64'b0001000000100000010000000101000001000000000000010000000000001000;
//				GR[2048:2111] <= 64'b0001000000100000010000000110000001000000000000010000000000001000;
//				GR[2112:2175] <= 64'b0001000000100000010000000101000001000000000000010000000000001000;
//				GR[2176:2239] <= 64'b0001000000100000010000000100100001000000000000010000000000001000;
//				GR[2240:2303] <= 64'b0001000000100000010000000100010001000000000000010000000000001000;
//				GR[2304:2367] <= 64'b0001000000100000010000000100001001000000000000010000000000001000;
//				GR[2368:2431] <= 64'b0001000000100000010000000100000101000000000000010000000000001000;
//				GR[2432:2495] <= 64'b0001000000100000010000000100000011000000000000010000000000001000;
//				GR[2496:2559] <= 64'b0001000000100000010000000100000101000000000000010000000000001000;
//				GR[2560:2623] <= 64'b0001000000100000010000000100001001000000000000010000000000001000;
//				GR[2624:2687] <= 64'b0001000000100000010000000100010001000001000000010000100000001000;
//				GR[2688:2751] <= 64'b0001000000100000010000000100100001000001000000010000100000001000;
//				GR[2752:2815] <= 64'b0001000000100000010000000101000001000001000000010000100000001000;
//				GR[2816:2879] <= 64'b0001000000100000010000000110000001000001000000010000100000001000;
//				GR[2880:2943] <= 64'b0001000000100000010000000111111111000001111111110000111111111000;
//				GR[2944:3007] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3008:3071] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3072:3135] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3136:3199] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
//				GR[3584:3647] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
//				GR[3648:3711] <= 64'b1110111011101110111011101110111011101110111011101110111011101110;
//				GR[3712:3775] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3776:3839] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3840:3903] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3904:3967] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[3968:4031] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//				GR[4032:4095] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
//			end
//		end
//	end
	
//	always @(state) begin
//		if(state==2'b01) begin
//			if(tmp_score_unit==9) begin
//				tmp_score_tens <= (tmp_score_tens+1);
//				tmp_score_unit <= 0;
//			end
//			else begin
//				tmp_score_unit <= (tmp_score_unit+1);
//			end
//		end
//		else begin
//		end
//	end
	
	// Control the output game view(Right)
//	always @(state) begin
//		case(state)
//			2'b01: begin
//				
//			end
//			2'b10: begin
//				
//			end
//			default: begin
//				
//			end
//		endcase
//	end
	
	// Control the output game view(Left)
	always @(posedge clk_1s or negedge reset) begin
		if(!reset) begin // Reset state, so the graph only has a rectangle at the middle of the LCD
			GL[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[  64: 127] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 128: 191] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 192: 255] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 256: 319] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 320: 383] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[ 832: 895] <= 64'b0011111111111111111111111111111111111111111111111111111111111100;
			GL[ 896: 959] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[ 960:1023] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1024:1087] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1088:1151] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1152:1215] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1216:1279] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1280:1343] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1344:1407] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1408:1471] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1472:1535] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1536:1599] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1600:1663] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1664:1727] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1728:1791] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1792:1855] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1856:1919] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1920:1983] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[1984:2047] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2048:2111] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2112:2175] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2176:2239] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2240:2303] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2304:2367] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2368:2431] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2432:2495] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2496:2559] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2560:2623] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2624:2687] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2688:2751] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2752:2815] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2816:2879] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2880:2943] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[2944:3007] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[3008:3071] <= 64'b0010000000000000000000000000000000000000000000000000000000000100;
			GL[3072:3135] <= 64'b0011111111111111111111111111111111111111111111111111111111111100;
			GL[3136:3199] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3584:3647] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3648:3711] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3712:3775] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			GL[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
		end
		else begin
			case(Melody)
				4'b0000: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000110000000000000000110000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000100000000000000000010000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000110000000000000000110000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b00001: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111100000000000000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000111111111111111111111111100000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b0010: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000111111111111111111000000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000111111111111111111000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000100000000000000000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000111111111111111111000000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b0011: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000111111111111111111000000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000111111111111111111000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000000000000000000001000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000111111111111111111000000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b0100: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000010000000100000000000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000000000000100000000000000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b0101: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b0110: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b0111: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1000: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1001: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000000000000000000000100000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1010: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1011: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111110000000000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000001000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000100000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000010000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000010000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000100000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000000001000000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000011111111111110000000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000001000000000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000100000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000010000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000000010000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000000100000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000000001000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111111110000000000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1100: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111000000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1101: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111110000000000000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000001000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000100000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000010000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000001000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000100000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000010000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000000100000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000001000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000010000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000100000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000001000000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000010000000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000100000000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000001000000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111110000000000000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1110: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4'b1111: begin
					GL[0:63]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[64:127]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[128:191]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[192:255]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[256:319]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[320:383]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[384:447]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[448:511]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[512:575]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[576:639]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[640:703]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[704:767]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[768:831]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[832:895]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[896:959]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[960:1023]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1024:1087]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[1088:1151]<=64'b0010000000000000000000011111111111111111100000000000000000000100;
					GL[1152:1215]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1216:1279]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1280:1343]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1344:1407]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1408:1471]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1472:1535]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1536:1599]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1600:1663]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1664:1727]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1728:1791]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1792:1855]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1856:1919]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[1920:1983]<=64'b0010000000000000000000011111111111111100000000000000000000000100;
					GL[1984:2047]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2048:2111]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2112:2175]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2176:2239]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2240:2303]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2304:2367]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2368:2431]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2432:2495]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2496:2559]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2560:2623]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2624:2687]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2688:2751]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2752:2815]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2816:2879]<=64'b0010000000000000000000010000000000000000000000000000000000000100;
					GL[2880:2943]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[2944:3007]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3008:3071]<=64'b0010000000000000000000000000000000000000000000000000000000000100;
					GL[3072:3135]<=64'b0011111111111111111111111111111111111111111111111111111111111100;
					GL[3136:3199]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3200:3263]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3264:3327]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3328:3391]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3392:3455]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3456:3519]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3520:3583]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3584:3647]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3648:3711]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3712:3775]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3776:3839]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3840:3903]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3904:3967]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[3968:4031]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
					GL[4032:4095]<=64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
			endcase
		end
	end
	
//	assign score_tens = tmp_score_tens;
//	assign score_unit = tmp_score_unit;
	
endmodule
