`timescale 1ns / 1ps
module LCD_DISPLAY_CTRL(LEFT_GRAPH, RIGHT_GRAPH, GL, GR, LCD_state, Mode_state, reset, clk_LCD, clk_10Hz, clk_100Hz);

	input reset, clk_LCD, clk_10Hz, clk_100Hz;
	input LCD_state;
	input [1:0] Mode_state;
//	input [3:0] KEY_IN;
	input [0:4095] GL;
	input [0:4095] GR;
	
	output reg [0:4095] LEFT_GRAPH;
	output reg [0:4095] RIGHT_GRAPH;
	
	reg [0:4095] ML;
	reg [0:4095] MR;
	reg [0:4095] GGR;
	reg [2:0] counter = 0;
	reg [2:0] count = 0;
	reg [3:0] display = 0;
//	reg LCD_state;
//	reg [1:0] Mode_state;
	
	//Menu_Display menu_display(ML, MR, Mode_state, reset, clk);
	
	// Decide which graph to show, the Game View or the Menu View
//	always @(posedge clk_LCD or negedge reset) begin
//		if(!reset) begin
//			LEFT_GRAPH <= ML;
//			RIGHT_GRAPH <= MR;
//		end
//		else begin
//			if(LCD_state==0) begin
//				LEFT_GRAPH <= ML;
//				RIGHT_GRAPH <= MR;
//			end
//			else begin
//				LEFT_GRAPH <= GL;
//				RIGHT_GRAPH <= GR;
//			end
//		end
//	end
	
	always @(*) begin
		if(LCD_state==0) begin
			LEFT_GRAPH <= ML;
			RIGHT_GRAPH <= MR;
		end
		else begin
			LEFT_GRAPH <= GL;
			RIGHT_GRAPH <= GGR;
		end
	end
	
	
	// Control of the Menu View(Left)
	always @(posedge clk_10Hz or negedge reset) begin
		if(!reset) begin
			ML[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[  64: 127] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 128: 191] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 192: 255] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 256: 319] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 320: 383] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[ 640: 703] <= 64'b0000000000000011111111111111111111111111111100000000000000000000;
			ML[ 704: 767] <= 64'b0000000000111110000000100001100000000000000010000000000000000000;
			ML[ 768: 831] <= 64'b0000000000100000000011100011000000000000000001000000000000000000;
			ML[ 832: 895] <= 64'b0000000111100000000110000110000000000000000001110000000000000000;
			ML[ 896: 959] <= 64'b0000001110000000001100000100000000000000000000011000000000000000;
			ML[ 960:1023] <= 64'b0000110100000000011000001000000000000000000000000100000000000000;
			ML[1024:1087] <= 64'b0001101100000000010000010000000000000000000000000110000000000000;
			ML[1088:1151] <= 64'b0011001000000000110000010000000000000000000000000010000000000000;
			ML[1152:1215] <= 64'b0010011000000000110000110000000111000000011100000011000000000000;
			ML[1216:1279] <= 64'b0110010000000001100000100000001111100000111110000011000000000000;
			ML[1280:1343] <= 64'b0100010000000001000000100000011111110001111111000001100000000000;
			ML[1344:1407] <= 64'b0100010000000001000000100000011111110001111111000001100000000000;
			ML[1408:1471] <= 64'b0100010000000001000000100000011110010001111001000000100000000000;
			ML[1472:1535] <= 64'b0100010000000001000000100000011110010001111001000000100000000000;
			ML[1536:1599] <= 64'b1000010000000001000000100000001111110000111111000000100000000000;
			ML[1600:1663] <= 64'b1000010000000001000000100000000000000000000000000000100000000000;
			ML[1664:1727] <= 64'b1000010000000001000000100000100000000100000000100000100000000000;
			ML[1728:1791] <= 64'b1000010000000001000000100000111000000100000000100000100000000000;
			ML[1792:1855] <= 64'b1000010000000001000000100000011100001110000001100000100000000000;
			ML[1856:1919] <= 64'b1000010000000001000000100000000110011011000011000000100000000000;
			ML[1920:1983] <= 64'b1000010000000001000000100000000011110001111110000000100000000000;
			ML[1984:2047] <= 64'b0100001000000001000000100000000010000000000100000001100000000000;
			ML[2048:2111] <= 64'b0100001100000001000000110000000010000000000100000001000000000000;
			ML[2112:2175] <= 64'b0010000110000001100000111000000010000000000100000011000000000000;
			ML[2176:2239] <= 64'b0011000010000000110000011000000011000000001100000011000000000000;
			ML[2240:2303] <= 64'b0001000011000000011100001100000001100000011000000010000000000000;
			ML[2304:2367] <= 64'b0001100001000000000100000110000000111111110000000100000000000000;
			ML[2368:2431] <= 64'b0000100001100000000111000011000000000000000000001100000000000000;
			ML[2432:2495] <= 64'b0000011000100000000001100001100000000000000000011000000000000000;
			ML[2496:2559] <= 64'b0000001110100000000000110000110000000000000000110000000000000000;
			ML[2560:2623] <= 64'b0000000011011000000000001000001000000000000000100000000000000000;
			ML[2624:2687] <= 64'b0000000001001000000000001100001000000000000000100000000000000000;
			ML[2688:2751] <= 64'b0000000001111111111111111111111100000000000011100000000000000000;
			ML[2752:2815] <= 64'b0000000000000000000000000000011111111111111110000000000000000000;
			ML[2816:2879] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[2880:2943] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[2944:3007] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3008:3071] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3072:3135] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3136:3199] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3584:3647] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3648:3711] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3712:3775] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			ML[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
		end
		else begin
			case(counter)
				0: begin
					ML[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[  64: 127] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 128: 191] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 192: 255] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 256: 319] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 320: 383] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 640: 703] <= 64'b0000000000000011111111111111111111111111111100000000000000000000;
					ML[ 704: 767] <= 64'b0000000000111110000000110000011000000000000010000000000000011110;
					ML[ 768: 831] <= 64'b0000000000100000000011000000110000000000000001000000000000110011;
					ML[ 832: 895] <= 64'b0000000111100000000110000011100000000000000001110000000001100001;
					ML[ 896: 959] <= 64'b0000001110000000001100000110000000000000000000011000000001000001;
					ML[ 960:1023] <= 64'b0000110100000000011000001100000000000000000000000100000001000001;
					ML[1024:1087] <= 64'b0001101100000000010000001000000000000000000000000110000001000001;
					ML[1088:1151] <= 64'b0011001000000000100000011000000000000000000000000010000001000001;
					ML[1152:1215] <= 64'b0010011000000000100000010000000111000000011100000011000011000001;
					ML[1216:1279] <= 64'b0110010000000000100000010000001111100000111110000011100110000001;
					ML[1280:1343] <= 64'b0100010000000000100000010000011111110001111111000001101100000001;
					ML[1344:1407] <= 64'b0100010000000001100000110000011111110001111111000001111000000001;
					ML[1408:1471] <= 64'b0100010000000001000000100000011110010001111001000000100000000001;
					ML[1472:1535] <= 64'b0100010000000001000000100000011110010001111001000000100000000011;
					ML[1536:1599] <= 64'b1000010000000001000000100000001111110000111111000000100000000100;
					ML[1600:1663] <= 64'b1000010000000001000000100000000000000000000000000000100000011000;
					ML[1664:1727] <= 64'b1000010000000001000000100000100000000100000000100000100001110000;
					ML[1728:1791] <= 64'b1000010000000001000000100000111000000100000000100000100011000000;
					ML[1792:1855] <= 64'b1000010000000001000000100000011100001110000001100000100010000000;
					ML[1856:1919] <= 64'b1000010000000001000000100000000110011011000011000000101110000000;
					ML[1920:1983] <= 64'b1000010000000000100000100000000011110001111110000000111000000000;
					ML[1984:2047] <= 64'b0100001000000000100000110000000010000000000100000001100000000000;
					ML[2048:2111] <= 64'b0100001100000000110000010000000010000000000100000001000000000000;
					ML[2112:2175] <= 64'b0010000110000000011000011000000010000000000100000011000000000000;
					ML[2176:2239] <= 64'b0011000010000000001100001000000011000000001100000011000000000000;
					ML[2240:2303] <= 64'b0001000011000000000100001100000001100000011000000010000000000000;
					ML[2304:2367] <= 64'b0001100001000000000110000110000000111111110000000100000000000000;
					ML[2368:2431] <= 64'b0000100001100000000011000011000000000000000000001100000000000000;
					ML[2432:2495] <= 64'b0000011000100000000001100001100000000000000000011000000000000000;
					ML[2496:2559] <= 64'b0000001110010000000000110000110000000000000000110000000000000000;
					ML[2560:2623] <= 64'b0000000011001100000000001000001000000000000000100000000000000000;
					ML[2624:2687] <= 64'b0000000001000110000000001100001100000000000001100000000000000000;
					ML[2688:2751] <= 64'b0000000001111111111111111100000011000000000111000000000000000000;
					ML[2752:2815] <= 64'b0000000000000000000000000100000001111111111000000000000000000000;
					ML[2816:2879] <= 64'b0000000000000000000000000111000000110000000000000000000000000000;
					ML[2880:2943] <= 64'b0000000000000000000000000001000000011000000000000000000000000000;
					ML[2944:3007] <= 64'b0000000000000000000000000001100000001100000011110000000000000000;
					ML[3008:3071] <= 64'b0000000000000000000000000000110000000110000110011100000000000000;
					ML[3072:3135] <= 64'b0000000000000000000000000000011000000011001100000110000000000000;
					ML[3136:3199] <= 64'b0000000000000000000000000000001100000001101000000010000000000000;
					ML[3200:3263] <= 64'b0000000000000000000000000000000110000000111000000010000000000000;
					ML[3264:3327] <= 64'b0000000000000000000000000000000011000000000000000010000000000000;
					ML[3328:3391] <= 64'b0000000000000000000000000000000001100000000000000110000000000000;
					ML[3392:3455] <= 64'b0000000000000000000000000000000000011000000000000100000000000000;
					ML[3456:3519] <= 64'b0000000000000000000000000000000000000111110000001100000000000000;
					ML[3520:3583] <= 64'b0000000000000000000000000000000000000011111110111000000000000000;
					ML[3584:3647] <= 64'b0000000000000000000000000000000000000000000011100000000000000000;
					ML[3648:3711] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3712:3775] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				1: begin
					ML[   0:  63] <= 64'b0000000000000000000000000000000000000000000000001111000000000000;
					ML[  64: 127] <= 64'b0000000000000000000000000000000000000000000000110001111000000000;
					ML[ 128: 191] <= 64'b0000000000000000000000000000000000000000000001100000001110000000;
					ML[ 192: 255] <= 64'b0000000000000000000000000000000000000000000001000000000011000000;
					ML[ 256: 319] <= 64'b0000000000000000000000000000000000000000000001000000000001100000;
					ML[ 320: 383] <= 64'b0000000000000000000000000000000000000000000001100000000000100000;
					ML[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000011000000000100000;
					ML[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000001100000000100000;
					ML[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000100000000100000;
					ML[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000100000000100000;
					ML[ 640: 703] <= 64'b0000000000000011111111111111111111111111111100000100000000100000;
					ML[ 704: 767] <= 64'b0000000000111110000000110000011000000000000010000100000000100000;
					ML[ 768: 831] <= 64'b0000000000100000000011000000110000000000000001001100000000100000;
					ML[ 832: 895] <= 64'b0000000111100000000110000011100000000000000001111000000001100000;
					ML[ 896: 959] <= 64'b0000001110000000001100000110000000000000000000011000000011000000;
					ML[ 960:1023] <= 64'b0000110100000000011000001100000000000000000000000100000110000000;
					ML[1024:1087] <= 64'b0001101100000000010000001000000000000000000000000110001100000000;
					ML[1088:1151] <= 64'b0011001000000000100000011000000000000000000000000010111000000000;
					ML[1152:1215] <= 64'b0010011000000000100000010000000111000000011100000011100000000000;
					ML[1216:1279] <= 64'b0110010000000000100000010000001111100000111110000011100000000000;
					ML[1280:1343] <= 64'b0100010000000000100000010000011111110001111111000001100000000000;
					ML[1344:1407] <= 64'b0100010000000001100000110000011111110001111111000001100000000000;
					ML[1408:1471] <= 64'b0100010000000001000000100000011110010001111001000000100000000000;
					ML[1472:1535] <= 64'b0100010000000001000000100000011110010001111001000000100000000000;
					ML[1536:1599] <= 64'b1000010000000001000000100000001111110000111111000000100000000000;
					ML[1600:1663] <= 64'b1000010000000001000000100000000000000000000000000000100000000000;
					ML[1664:1727] <= 64'b1000010000000001000000100000100000000100000000100000100000000000;
					ML[1728:1791] <= 64'b1000010000000001000000100000111000000100000000100000100000000000;
					ML[1792:1855] <= 64'b1000010000000001000000100000011100001110000001100000100000000000;
					ML[1856:1919] <= 64'b1000010000000001000000100000000110011011000011000000100000000000;
					ML[1920:1983] <= 64'b1000010000000000100000100000000011110001111110000000100000000000;
					ML[1984:2047] <= 64'b0100001000000000100000110000000010000000000100000001100000000000;
					ML[2048:2111] <= 64'b0100001100000000110000010000000010000000000100000001000000000000;
					ML[2112:2175] <= 64'b0010000110000000011000011000000010000000000100000011000000000000;
					ML[2176:2239] <= 64'b0011000010000000001100001000000011000000001100000011000000000000;
					ML[2240:2303] <= 64'b0001000011000000000100001100000001100000011000000010000000000000;
					ML[2304:2367] <= 64'b0001100001000000000110000110000000111111110000000100000000000000;
					ML[2368:2431] <= 64'b0000100001100000000011000011000000000000000000001100000000000000;
					ML[2432:2495] <= 64'b0000011000100000000001100001100000000000000000011000000000000000;
					ML[2496:2559] <= 64'b0000001110010000000000110000110000000000000000110000000000000000;
					ML[2560:2623] <= 64'b0000000011001100000000001000001000000000000000100000000000000000;
					ML[2624:2687] <= 64'b0000000001000110000000001100001100000000000001100000000000000000;
					ML[2688:2751] <= 64'b0000000001111111111111111100000011000000000111000000000000000000;
					ML[2752:2815] <= 64'b0000000000000000000000000110000001111111111000000000000011111000;
					ML[2816:2879] <= 64'b0000000000000000000000000001110000011111110000000000001100001100;
					ML[2880:2943] <= 64'b0000000000000000000000000000011100000000011111000000011000000110;
					ML[2944:3007] <= 64'b0000000000000000000000000000000111100000000001110000110000000010;
					ML[3008:3071] <= 64'b0000000000000000000000000000000000111000000000011111100000000010;
					ML[3072:3135] <= 64'b0000000000000000000000000000000000001100000000000000000000000001;
					ML[3136:3199] <= 64'b0000000000000000000000000000000000000111000000000000000000000001;
					ML[3200:3263] <= 64'b0000000000000000000000000000000000000000111000000000000000000011;
					ML[3264:3327] <= 64'b0000000000000000000000000000000000000000001111000000000000000110;
					ML[3328:3391] <= 64'b0000000000000000000000000000000000000000000000111111000000011100;
					ML[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000001111111110000;
					ML[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3584:3647] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3648:3711] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3712:3775] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				2: begin
					ML[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[  64: 127] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 128: 191] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 192: 255] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 256: 319] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 320: 383] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 448: 511] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 512: 575] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 576: 639] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[ 640: 703] <= 64'b0000000000000011111111111111111111111111111100000000000000000000;
					ML[ 704: 767] <= 64'b0000000000111110000000100001100000000000000010000000000000000000;
					ML[ 768: 831] <= 64'b0000000000100000000011100011000000000000000001000000000000000000;
					ML[ 832: 895] <= 64'b0000000111100000000110000110000000000000000001110000000000000000;
					ML[ 896: 959] <= 64'b0000001110000000001100000100000000000000000000011000000000000000;
					ML[ 960:1023] <= 64'b0000110100000000011000001000000000000000000000000100000000000000;
					ML[1024:1087] <= 64'b0001101100000000010000010000000000000000000000000110000000000000;
					ML[1088:1151] <= 64'b0011001000000000110000010000000000000000000000000010000011111110;
					ML[1152:1215] <= 64'b0010011000000000110000110000000111000000011100000011000110000011;
					ML[1216:1279] <= 64'b0110010000000001100000100000001111100000111110000011001100000001;
					ML[1280:1343] <= 64'b0100010000000001000000100000011111110001111111000001101000000001;
					ML[1344:1407] <= 64'b0100010000000001000000100000011111110001111111000001101000000001;
					ML[1408:1471] <= 64'b0100010000000001000000100000011110010001111001000000101000000001;
					ML[1472:1535] <= 64'b0100010000000001000000100000011110010001111001000000101100000001;
					ML[1536:1599] <= 64'b1000010000000001000000100000001111110000111111000000100100000011;
					ML[1600:1663] <= 64'b1000010000000001000000100000000000000000000000000000100100000010;
					ML[1664:1727] <= 64'b1000010000000001000000100000100000000100000000100000101100000010;
					ML[1728:1791] <= 64'b1000010000000001000000100000111000000100000000100000111000000110;
					ML[1792:1855] <= 64'b1000010000000001000000100000011100001110000001100000110000000100;
					ML[1856:1919] <= 64'b1000010000000001000000100000000110011011000011000001100000001100;
					ML[1920:1983] <= 64'b1000010000000001000000100000000011110001111110000011000000011000;
					ML[1984:2047] <= 64'b0100001000000001000000100000000010000000000100000110000000110000;
					ML[2048:2111] <= 64'b0100001100000001000000110000000010000000000100001100000001100000;
					ML[2112:2175] <= 64'b0010000110000001100000111000000010000000000100011000000011000000;
					ML[2176:2239] <= 64'b0011000010000000110000011000000011000000001100110000000110000000;
					ML[2240:2303] <= 64'b0001000011000000011100001100000001100000011111100000011000000000;
					ML[2304:2367] <= 64'b0001100001000000000100000110000000111111111000000001110000000000;
					ML[2368:2431] <= 64'b0000100001100000000111000011000000000001100000000111000001111110;
					ML[2432:2495] <= 64'b0000011000100000000001100001100000001110000000001110000001000011;
					ML[2496:2559] <= 64'b0000001110100000000000110000110000111000000000011100000011000001;
					ML[2560:2623] <= 64'b0000000011011000000000001000001111100000000000110110000011000001;
					ML[2624:2687] <= 64'b0000000001001000000000001100001100000000000001100011100111000001;
					ML[2688:2751] <= 64'b0000000001111111111111111110000110000000000011100000111100000001;
					ML[2752:2815] <= 64'b0000000000000000000000000011111111111111111111000000000000000011;
					ML[2816:2879] <= 64'b0000000000000000000000000000000000000000000000110000000000000110;
					ML[2880:2943] <= 64'b0000000000000000000000000000000000000000000000011000000000000110;
					ML[2944:3007] <= 64'b0000000000000000000000000000000000000000000000001110000000000100;
					ML[3008:3071] <= 64'b0000000000000000000000000000000000000000000000000011110000011100;
					ML[3072:3135] <= 64'b0000000000000000000000000000000000000000000000000000001111110000;
					ML[3136:3199] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3584:3647] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3648:3711] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3712:3775] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				3: begin
					ML[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[  64: 127] <= 64'b0000000000000000001111111100000000000000000000000000000000000000;
					ML[ 128: 191] <= 64'b0000000000000000110000000011110000000000000000000000000000000000;
					ML[ 192: 255] <= 64'b0000000000000001100000000000011000000000000000000000000000000000;
					ML[ 256: 319] <= 64'b0000000000000001000000000000001000000000000000000000000000000000;
					ML[ 320: 383] <= 64'b0000000000000001000000000000001000000000000000000000000000000000;
					ML[ 384: 447] <= 64'b0000000000000001100000000000001000000000000000000000000000000000;
					ML[ 448: 511] <= 64'b0000000000000000111100000000001000000000000000000000000000000000;
					ML[ 512: 575] <= 64'b0000000000000000000111100000001000000000000000000000000000000000;
					ML[ 576: 639] <= 64'b0000000000000000000001100000011000000000000000000000000000000000;
					ML[ 640: 703] <= 64'b0000000000000011111111100000011111111111111100000000000000000000;
					ML[ 704: 767] <= 64'b0000000000111110000000100000011000000000000010000000000000000000;
					ML[ 768: 831] <= 64'b0000000000100000000011100000010000000000000001000000000000000000;
					ML[ 832: 895] <= 64'b0000000111100000000110100000010000000000000001110000000000000000;
					ML[ 896: 959] <= 64'b0000001110000000001100100000110000000000000000011000000000000000;
					ML[ 960:1023] <= 64'b0000110100000000011000100000100000000000000000000100000000000000;
					ML[1024:1087] <= 64'b0001101100000000010000100000100000000000000000000110000000000000;
					ML[1088:1151] <= 64'b0011001000000000100000100000100000000000000000000010000000000000;
					ML[1152:1215] <= 64'b0010011000000000100000100001100111000000011100000011000000000000;
					ML[1216:1279] <= 64'b0110010000000000100000100001001111100000111110000011000000000000;
					ML[1280:1343] <= 64'b0100010000000000100001000001011111110001111111000001100000000000;
					ML[1344:1407] <= 64'b0100010000000001100001000011011111110001111111000001100000000000;
					ML[1408:1471] <= 64'b0100010000000001000010000010011110010001111001000000100000000000;
					ML[1472:1535] <= 64'b0100010000000001000110000010011110010001111001000000100000000000;
					ML[1536:1599] <= 64'b1000010000000001000100000100001111110000111111000000100000000000;
					ML[1600:1663] <= 64'b1000010000000001001000000100000000000000000000000000100000000000;
					ML[1664:1727] <= 64'b1000010000000001001000001100100000000100000000100000100000000000;
					ML[1728:1791] <= 64'b1000010000000001011000001000111000000100000000100000100000000000;
					ML[1792:1855] <= 64'b1000010000000001010000011000011100001110000001100000100000000000;
					ML[1856:1919] <= 64'b1000010000000001010000010000000110011011000011000000100000000000;
					ML[1920:1983] <= 64'b1000010000000001110000010000000011110001111110000000100000000000;
					ML[1984:2047] <= 64'b0100001000000001000000010000000010000000000100000001100000000000;
					ML[2048:2111] <= 64'b0100001100000001000000110000000010000000000100000001000000000000;
					ML[2112:2175] <= 64'b0010000110000001000001011000000010000000000100000011000000000000;
					ML[2176:2239] <= 64'b0011000010000011000001001000000011000000001100000011000000000000;
					ML[2240:2303] <= 64'b0001000011000110000011001100000001100000011000000010000000000000;
					ML[2304:2367] <= 64'b0001100001000100000010000110000000111111110000000100000000000000;
					ML[2368:2431] <= 64'b0000100001101000000111000011000000000000000000001100000000000000;
					ML[2432:2495] <= 64'b0000011000110000001101100001100000000000000000011000000000000000;
					ML[2496:2559] <= 64'b0000001110010000001100110000110000000000000000110000000000000000;
					ML[2560:2623] <= 64'b0000000011010000011000001000001000000000000011100000000000000000;
					ML[2624:2687] <= 64'b0000000001011110110000001100001000000000000011000000000000000000;
					ML[2688:2751] <= 64'b0000000001111111111111111111111111000000000011100000001111100000;
					ML[2752:2815] <= 64'b0000000000000000000000000000011111111111111111110000011000100000;
					ML[2816:2879] <= 64'b0000000000000000000000000000000000000011000000011000110000010000;
					ML[2880:2943] <= 64'b0000000000000000000000000000000000000001000000000110100000011000;
					ML[2944:3007] <= 64'b0000000000000000000000000000000000000001100000000011100000001000;
					ML[3008:3071] <= 64'b0000000000000000000000000000000000000000110000000001100000001000;
					ML[3072:3135] <= 64'b0000000000000000000000000000000000000000011100000000000000001000;
					ML[3136:3199] <= 64'b0000000000000000000000000000000000000000000110000000000000011000;
					ML[3200:3263] <= 64'b0000000000000000000000000000000000000000000011000000000000110000;
					ML[3264:3327] <= 64'b0000000000000000000000000000000000000000000000110000000001100000;
					ML[3328:3391] <= 64'b0000000000000000000000000000000000000000000000011000000110000000;
					ML[3392:3455] <= 64'b0000000000000000000000000000000000000000000000000111111000000000;
					ML[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3520:3583] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3584:3647] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3648:3711] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3712:3775] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					ML[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
			endcase
			if(counter==3'b100)
				counter <= 3'b000;
			else
				counter <= (counter+1);
		end
	end
	
	// Control of the Menu View(Right)
	always @(posedge clk_LCD or negedge reset) begin
		if(!reset) begin
			MR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[  64: 127] <= 64'b0011111001111000100010010011110000000000000111110001111000111100;
			MR[ 128: 191] <= 64'b0000100000001000000010100010010000000000000001000000001000100100;
			MR[ 192: 255] <= 64'b0000100001111000100011000010010000000000000001000001111000111100;
			MR[ 256: 319] <= 64'b0000100001001000100010100010010000000000000001000001001000100000;
			MR[ 320: 383] <= 64'b0000100001111000100010010011110000000000000001000001111000100000;
			MR[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[ 448: 511] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
			MR[ 512: 575] <= 64'b1010101010101010101010101010101010101010101010101010101010101010;
			MR[ 576: 639] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
			MR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[ 832: 895] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
			MR[ 896: 959] <= 64'b0000000000000000100000001000100010001000100010000000000000000000;
			MR[ 960:1023] <= 64'b0000000000000000100000001000100010000000100010000000000000000000;
			MR[1024:1087] <= 64'b0000000000000000111110001111100011111000111110000000000000000000;
			MR[1088:1151] <= 64'b0000000000000000100000001000100000001000001000000000000000000000;
			MR[1152:1215] <= 64'b0000000000000000100000001000100010001000001000000000000000000000;
			MR[1216:1279] <= 64'b0000000000000000111110001000100011111000001000000000000000000000;
			MR[1280:1343] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1344:1407] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1408:1471] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1472:1535] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1536:1599] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1600:1663] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1664:1727] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1728:1791] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[1792:1855] <= 64'b0000000000111110001111100011111000111110001111100010000000000000;
			MR[1856:1919] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
			MR[1920:1983] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
			MR[1984:2047] <= 64'b0000000000100010001000100010000000101010001111100010000000000000;
			MR[2048:2111] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
			MR[2112:2175] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
			MR[2176:2239] <= 64'b0000000000100010001111100010000000101010001111100011111000000000;
			MR[2240:2303] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2304:2367] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2368:2431] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2432:2495] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2496:2559] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2560:2623] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2624:2687] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2688:2751] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[2752:2815] <= 64'b0000000000000000100010001111100011111000111000000000000000000000;
			MR[2816:2879] <= 64'b0000000000000000100010001000100010001000101100000000000000000000;
			MR[2880:2943] <= 64'b0000000000000000100010001000100010001000100110000000000000000000;
			MR[2944:3007] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
			MR[3008:3071] <= 64'b0000000000000000100010001000100011100000100110000000000000000000;
			MR[3072:3135] <= 64'b0000000000000000100010001000100010110000101100000000000000000000;
			MR[3136:3199] <= 64'b0000000000000000100010001000100010011000111000000000000000000000;
			MR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[3392:3455] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
			MR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			MR[3520:3583] <= 64'b0111000000000000001000000000100000000000000000011110001111011110;
			MR[3584:3647] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
			MR[3648:3711] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
			MR[3712:3775] <= 64'b0111010101011100001010001011101110100010111000011110101000010010;
			MR[3776:3839] <= 64'b0101000101010100001111100010101010101010101000000010001011010010;
			MR[3840:3903] <= 64'b0101010111011100000010001011101110111110101000000010101001010010;
			MR[3904:3967] <= 64'b0111000000010000000010000000000000000000000000011110001111011110;
			MR[3968:4031] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
			MR[4032:4095] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
		end
		else begin
			case(Mode_state)
				1: begin
					MR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[  64: 127] <= 64'b0011111001111000100010010011110000000000000111110001111000111100;
					MR[ 128: 191] <= 64'b0000100000001000000010100010010000000000000001000000001000100100;
					MR[ 192: 255] <= 64'b0000100001111000100011000010010000000000000001000001111000111100;
					MR[ 256: 319] <= 64'b0000100001001000100010100010010000000000000001000001001000100000;
					MR[ 320: 383] <= 64'b0000100001111000100010010011110000000000000001000001111000100000;
					MR[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[ 448: 511] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
					MR[ 512: 575] <= 64'b1010101010101010101010101010101010101010101010101010101010101010;
					MR[ 576: 639] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
					MR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[ 832: 895] <= 64'b0000010100000000111110001111100011111000100010000000000010100000;
					MR[ 896: 959] <= 64'b0000101000000000100000001000100010001000100010000000000001010000;
					MR[ 960:1023] <= 64'b0001010000000000100000001000100010000000100010000000000000101000;
					MR[1024:1087] <= 64'b0001010000000000111110001111100011111000111110000000000000101000;
					MR[1088:1151] <= 64'b0001010000000000100000001000100000001000001000000000000000101000;
					MR[1152:1215] <= 64'b0000101000000000100000001000100010001000001000000000000001010000;
					MR[1216:1279] <= 64'b0000010100000000111110001000100011111000001000000000000010100000;
					MR[1280:1343] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1344:1407] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1408:1471] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1472:1535] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1536:1599] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1600:1663] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1664:1727] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1728:1791] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[1792:1855] <= 64'b0000000000111110001111100011111000111110001111100010000000000000;
					MR[1856:1919] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
					MR[1920:1983] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
					MR[1984:2047] <= 64'b0000000000100010001000100010000000101010001111100010000000000000;
					MR[2048:2111] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
					MR[2112:2175] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
					MR[2176:2239] <= 64'b0000000000100010001111100010000000101010001111100011111000000000;
					MR[2240:2303] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2304:2367] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2368:2431] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2432:2495] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2496:2559] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2560:2623] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2624:2687] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2688:2751] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[2752:2815] <= 64'b0000000000000000100010001111100011111000111000000000000000000000;
					MR[2816:2879] <= 64'b0000000000000000100010001000100010001000101100000000000000000000;
					MR[2880:2943] <= 64'b0000000000000000100010001000100010001000100110000000000000000000;
					MR[2944:3007] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
					MR[3008:3071] <= 64'b0000000000000000100010001000100011100000100110000000000000000000;
					MR[3072:3135] <= 64'b0000000000000000100010001000100010110000101100000000000000000000;
					MR[3136:3199] <= 64'b0000000000000000100010001000100010011000111000000000000000000000;
					MR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[3392:3455] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
					MR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					MR[3520:3583] <= 64'b0111000000000000001000000000100000000000000000011110001111011110;
					MR[3584:3647] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
					MR[3648:3711] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
					MR[3712:3775] <= 64'b0111010101011100001010001011101110100010111000011110101000010010;
					MR[3776:3839] <= 64'b0101000101010100001111100010101010101010101000000010001011010010;
					MR[3840:3903] <= 64'b0101010111011100000010001011101110111110101000000010101001010010;
					MR[3904:3967] <= 64'b0111000000010000000010000000000000000000000000011110001111011110;
					MR[3968:4031] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
					MR[4032:4095] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
				end
			2: begin
				MR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[  64: 127] <= 64'b0011111001111000100010010011110000000000000111110001111000111100;
				MR[ 128: 191] <= 64'b0000100000001000000010100010010000000000000001000000001000100100;
				MR[ 192: 255] <= 64'b0000100001111000100011000010010000000000000001000001111000111100;
				MR[ 256: 319] <= 64'b0000100001001000100010100010010000000000000001000001001000100000;
				MR[ 320: 383] <= 64'b0000100001111000100010010011110000000000000001000001111000100000;
				MR[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 448: 511] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
				MR[ 512: 575] <= 64'b1010101010101010101010101010101010101010101010101010101010101010;
				MR[ 576: 639] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
				MR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 832: 895] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
				MR[ 896: 959] <= 64'b0000000000000000100000001000100010001000100010000000000000000000;
				MR[ 960:1023] <= 64'b0000000000000000100000001000100010000000100010000000000000000000;
				MR[1024:1087] <= 64'b0000000000000000111110001111100011111000111110000000000000000000;
				MR[1088:1151] <= 64'b0000000000000000100000001000100000001000001000000000000000000000;
				MR[1152:1215] <= 64'b0000000000000000100000001000100010001000001000000000000000000000;
				MR[1216:1279] <= 64'b0000000000000000111110001000100011111000001000000000000000000000;
				MR[1280:1343] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1344:1407] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1408:1471] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1472:1535] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1536:1599] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1600:1663] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1664:1727] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1728:1791] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1792:1855] <= 64'b0000010100111110001111100011111000111110001111100010000010100000;
				MR[1856:1919] <= 64'b0000101000100010001000100010000000101010000000100010000001010000;
				MR[1920:1983] <= 64'b0001010000100010001000100010000000101010000000100010000000101000;
				MR[1984:2047] <= 64'b0001010000100010001000100010000000101010001111100010000000101000;
				MR[2048:2111] <= 64'b0001010000100010001000100010000000101010001000100010000000101000;
				MR[2112:2175] <= 64'b0000101000100010001000100010000000101010001000100010000001010000;
				MR[2176:2239] <= 64'b0000010100100010001111100010000000101010001111100011111010100000;
				MR[2240:2303] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2304:2367] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2368:2431] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2432:2495] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2496:2559] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2560:2623] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2624:2687] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2688:2751] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2752:2815] <= 64'b0000000000000000100010001111100011111000111000000000000000000000;
				MR[2816:2879] <= 64'b0000000000000000100010001000100010001000101100000000000000000000;
				MR[2880:2943] <= 64'b0000000000000000100010001000100010001000100110000000000000000000;
				MR[2944:3007] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
				MR[3008:3071] <= 64'b0000000000000000100010001000100011100000100110000000000000000000;
				MR[3072:3135] <= 64'b0000000000000000100010001000100010110000101100000000000000000000;
				MR[3136:3199] <= 64'b0000000000000000100010001000100010011000111000000000000000000000;
				MR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3392:3455] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
				MR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3520:3583] <= 64'b0111000000000000001000000000100000000000000000011110001111011110;
				MR[3584:3647] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
				MR[3648:3711] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
				MR[3712:3775] <= 64'b0111010101011100001010001011101110100010111000011110101000010010;
				MR[3776:3839] <= 64'b0101000101010100001111100010101010101010101000000010001011010010;
				MR[3840:3903] <= 64'b0101010111011100000010001011101110111110101000000010101001010010;
				MR[3904:3967] <= 64'b0111000000010000000010000000000000000000000000011110001111011110;
				MR[3968:4031] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
				MR[4032:4095] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
			end
			3: begin
				MR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[  64: 127] <= 64'b0011111001111000100010010011110000000000000111110001111000111100;
				MR[ 128: 191] <= 64'b0000100000001000000010100010010000000000000001000000001000100100;
				MR[ 192: 255] <= 64'b0000100001111000100011000010010000000000000001000001111000111100;
				MR[ 256: 319] <= 64'b0000100001001000100010100010010000000000000001000001001000100000;
				MR[ 320: 383] <= 64'b0000100001111000100010010011110000000000000001000001111000100000;
				MR[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 448: 511] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
				MR[ 512: 575] <= 64'b1010101010101010101010101010101010101010101010101010101010101010;
				MR[ 576: 639] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
				MR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 832: 895] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
				MR[ 896: 959] <= 64'b0000000000000000100000001000100010001000100010000000000000000000;
				MR[ 960:1023] <= 64'b0000000000000000100000001000100010000000100010000000000000000000;
				MR[1024:1087] <= 64'b0000000000000000111110001111100011111000111110000000000000000000;
				MR[1088:1151] <= 64'b0000000000000000100000001000100000001000001000000000000000000000;
				MR[1152:1215] <= 64'b0000000000000000100000001000100010001000001000000000000000000000;
				MR[1216:1279] <= 64'b0000000000000000111110001000100011111000001000000000000000000000;
				MR[1280:1343] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1344:1407] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1408:1471] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1472:1535] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1536:1599] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1600:1663] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1664:1727] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1728:1791] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1792:1855] <= 64'b0000000000111110001111100011111000111110001111100010000000000000;
				MR[1856:1919] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
				MR[1920:1983] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
				MR[1984:2047] <= 64'b0000000000100010001000100010000000101010001111100010000000000000;
				MR[2048:2111] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
				MR[2112:2175] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
				MR[2176:2239] <= 64'b0000000000100010001111100010000000101010001111100011111000000000;
				MR[2240:2303] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2304:2367] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2368:2431] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2432:2495] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2496:2559] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2560:2623] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2624:2687] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2688:2751] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2752:2815] <= 64'b0000010100000000100010001111100011111000111000000000000001010000;
				MR[2816:2879] <= 64'b0000101000000000100010001000100010001000101100000000000000101000;
				MR[2880:2943] <= 64'b0001010000000000100010001000100010001000100110000000000000010100;
				MR[2944:3007] <= 64'b0001010000000000111110001111100011111000100010000000000000010100;
				MR[3008:3071] <= 64'b0001010000000000100010001000100011100000100110000000000000010100;
				MR[3072:3135] <= 64'b0000101000000000100010001000100010110000101100000000000000101000;
				MR[3136:3199] <= 64'b0000010100000000100010001000100010011000111000000000000001010000;
				MR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3392:3455] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
				MR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3520:3583] <= 64'b0111000000000000001000000000100000000000000000011110001111011110;
				MR[3584:3647] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
				MR[3648:3711] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
				MR[3712:3775] <= 64'b0111010101011100001010001011101110100010111000011110101000010010;
				MR[3776:3839] <= 64'b0101000101010100001111100010101010101010101000000010001011010010;
				MR[3840:3903] <= 64'b0101010111011100000010001011101110111110101000000010101001010010;
				MR[3904:3967] <= 64'b0111000000010000000010000000000000000000000000011110001111011110;
				MR[3968:4031] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
				MR[4032:4095] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
			end
			default: begin
				MR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[  64: 127] <= 64'b0011111001111000100010010011110000000000000111110001111000111100;
				MR[ 128: 191] <= 64'b0000100000001000000010100010010000000000000001000000001000100100;
				MR[ 192: 255] <= 64'b0000100001111000100011000010010000000000000001000001111000111100;
				MR[ 256: 319] <= 64'b0000100001001000100010100010010000000000000001000001001000100000;
				MR[ 320: 383] <= 64'b0000100001111000100010010011110000000000000001000001111000100000;
				MR[ 384: 447] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 448: 511] <= 64'b0100010001000100010001000100010001000100010001000100010001000100;
				MR[ 512: 575] <= 64'b1010101010101010101010101010101010101010101010101010101010101010;
				MR[ 576: 639] <= 64'b0001000100010001000100010001000100010001000100010001000100010001;
				MR[ 640: 703] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 704: 767] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 768: 831] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[ 832: 895] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
				MR[ 896: 959] <= 64'b0000000000000000100000001000100010001000100010000000000000000000;
				MR[ 960:1023] <= 64'b0000000000000000100000001000100010000000100010000000000000000000;
				MR[1024:1087] <= 64'b0000000000000000111110001111100011111000111110000000000000000000;
				MR[1088:1151] <= 64'b0000000000000000100000001000100000001000001000000000000000000000;
				MR[1152:1215] <= 64'b0000000000000000100000001000100010001000001000000000000000000000;
				MR[1216:1279] <= 64'b0000000000000000111110001000100011111000001000000000000000000000;
				MR[1280:1343] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1344:1407] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1408:1471] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1472:1535] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1536:1599] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1600:1663] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1664:1727] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1728:1791] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[1792:1855] <= 64'b0000000000111110001111100011111000111110001111100010000000000000;
				MR[1856:1919] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
				MR[1920:1983] <= 64'b0000000000100010001000100010000000101010000000100010000000000000;
				MR[1984:2047] <= 64'b0000000000100010001000100010000000101010001111100010000000000000;
				MR[2048:2111] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
				MR[2112:2175] <= 64'b0000000000100010001000100010000000101010001000100010000000000000;
				MR[2176:2239] <= 64'b0000000000100010001111100010000000101010001111100011111000000000;
				MR[2240:2303] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2304:2367] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2368:2431] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2432:2495] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2496:2559] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2560:2623] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2624:2687] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2688:2751] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[2752:2815] <= 64'b0000000000000000100010001111100011111000111000000000000000000000;
				MR[2816:2879] <= 64'b0000000000000000100010001000100010001000101100000000000000000000;
				MR[2880:2943] <= 64'b0000000000000000100010001000100010001000100110000000000000000000;
				MR[2944:3007] <= 64'b0000000000000000111110001111100011111000100010000000000000000000;
				MR[3008:3071] <= 64'b0000000000000000100010001000100011100000100110000000000000000000;
				MR[3072:3135] <= 64'b0000000000000000100010001000100010110000101100000000000000000000;
				MR[3136:3199] <= 64'b0000000000000000100010001000100010011000111000000000000000000000;
				MR[3200:3263] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3264:3327] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3328:3391] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3392:3455] <= 64'b1111111111111111111111111111111111111111111111111111111111111111;
				MR[3456:3519] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				MR[3520:3583] <= 64'b0111000000000000001000000000100000000000000000011110001111011110;
				MR[3584:3647] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
				MR[3648:3711] <= 64'b0100000000000000001010000000100000000000000000010000001000010010;
				MR[3712:3775] <= 64'b0111010101011100001010001011101110100010111000011110101000010010;
				MR[3776:3839] <= 64'b0101000101010100001111100010101010101010101000000010001011010010;
				MR[3840:3903] <= 64'b0101010111011100000010001011101110111110101000000010101001010010;
				MR[3904:3967] <= 64'b0111000000010000000010000000000000000000000000011110001111011110;
				MR[3968:4031] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
				MR[4032:4095] <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
			end
			endcase
		end
	end
	
	always @(posedge clk_100Hz) begin
		if(display%7==0) begin
			case(count)
				0: begin
					GGR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[  64: 127] <= 64'b0000000000000000111111100000000000000000000000000000000000000000;
					GGR[ 128: 191] <= 64'b0000000000000011100000100000001111100000000000000000000000000000;
					GGR[ 192: 255] <= 64'b0000000000011111000001100011111000111000000000000000000000000000;
					GGR[ 256: 319] <= 64'b0000000000110000000011000000000000001110000000000000000000000000;
					GGR[ 320: 383] <= 64'b0000000001100000000110000000000000000001000000000000000000000000;
					GGR[ 384: 447] <= 64'b0000000001000000001100000000111111000000000000000000000000000000;
					GGR[ 448: 511] <= 64'b0000000011000000111000000000000000111000000000000000000000000000;
					GGR[ 512: 575] <= 64'b0000000010000001111000000000000000001000000000000000000000000000;
					GGR[ 576: 639] <= 64'b0000000010000001000000001111110000000000000000000000000000000000;
					GGR[ 640: 703] <= 64'b0000000011000001000000000000001000000000000000000000000000000000;
					GGR[ 704: 767] <= 64'b0000000001100001000000000000000000000000000000000000000000000000;
					GGR[ 768: 831] <= 64'b0000000000100000100001111111111111111111110000000000000000000000;
					GGR[ 832: 895] <= 64'b0000000000100000110011000000011100010000001111000000000000000000;
					GGR[ 896: 959] <= 64'b0000000000110000011110000000000100001100000000111100000000000000;
					GGR[ 960:1023] <= 64'b0000000000011000111100000000000110000100000000000111000000000000;
					GGR[1024:1087] <= 64'b0000000000001111100000000000000011000010000000000001100000000000;
					GGR[1088:1151] <= 64'b0000000000000110000000000000000001100001000000000000111000000000;
					GGR[1152:1215] <= 64'b0000000000011000000000000000000000100000100000000000011100000000;
					GGR[1216:1279] <= 64'b0000000000010000000000000000000000010000100000000000011110000000;
					GGR[1280:1343] <= 64'b0000000000100000000000000000000000011000100000000000001111000000;
					GGR[1344:1407] <= 64'b0000000000100000111100000001111000001000010000000000000101100000;
					GGR[1408:1471] <= 64'b0000000001000001111110000011111100000100010000000000000110110000;
					GGR[1472:1535] <= 64'b0000000001000011111111000011111110000100011000000000000010011000;
					GGR[1536:1599] <= 64'b0000000010000011111111000111111110000100001000000000000011001000;
					GGR[1600:1663] <= 64'b0000000010000010011111000110011110000100001000000000000001000100;
					GGR[1664:1727] <= 64'b0000000010000010011111000110011110000100001000000000000001000100;
					GGR[1728:1791] <= 64'b0000000010000011111111000011111110000100001000000000000001000110;
					GGR[1792:1855] <= 64'b0000000100000001111110000001111100000100001000000000000001000010;
					GGR[1856:1919] <= 64'b0000000100000000000000000000000000000100001000000000000001000010;
					GGR[1920:1983] <= 64'b0000000100000000000000000000000000000100001000000000000001000010;
					GGR[1984:2047] <= 64'b0000000100000110000000110000000001100100001000000000000001000010;
					GGR[2048:2111] <= 64'b0000000100000011000001111000000001000100001000000000000001000010;
					GGR[2112:2175] <= 64'b0000000100000001000011001000000011000100001000000000000001000010;
					GGR[2176:2239] <= 64'b0000000100000001100110001100000110001100001000000000000001000010;
					GGR[2240:2303] <= 64'b0000000010000001111100000111111110001000011000000000000001000010;
					GGR[2304:2367] <= 64'b0000000010000001000000000000000100001000110000000000000001000010;
					GGR[2368:2431] <= 64'b0000000011000001100000000000001100001000100000000000000001000010;
					GGR[2432:2495] <= 64'b0000000001000000100000000000011000011001100000000000000001000110;
					GGR[2496:2559] <= 64'b0000000001000000100000000000110000110001000000000000000011000100;
					GGR[2560:2623] <= 64'b0011111000100000010000000000100000100001000000000000000110001000;
					GGR[2624:2687] <= 64'b0110001100100000011000000011100001100011000000000000001100011000;
					GGR[2688:2751] <= 64'b1100000100010000001111111110000011000010000000000000001000010000;
					GGR[2752:2815] <= 64'b1000000110011000000000000000000010000110000000000000011001100000;
					GGR[2816:2879] <= 64'b1000000110001110000000000000001110001100000000000000010011000000;
					GGR[2880:2943] <= 64'b1000000110000111100000000000010000001000000000000000110110000000;
					GGR[2944:3007] <= 64'b1100000011111111111110000000110000011000000000000001111100000000;
					GGR[3008:3071] <= 64'b0100000000000000001111110001100000110000000000000011110000000000;
					GGR[3072:3135] <= 64'b0100000000000000000011111111100001100000000000000111000000000000;
					GGR[3136:3199] <= 64'b0011000000000000000000000000111111000000000000111100000000000000;
					GGR[3200:3263] <= 64'b0001110000000000000000000000001111111111111111110000000000000000;
					GGR[3264:3327] <= 64'b0100011100000000000000001111111100000000000000000000000000000000;
					GGR[3328:3391] <= 64'b0100000111110000011111111000000000000000000000000000000000000000;
					GGR[3392:3455] <= 64'b0110010000011111111110000000000000000000000000000000000000000000;
					GGR[3456:3519] <= 64'b0010010001000000000000000000000000000000000000000000000000000000;
					GGR[3520:3583] <= 64'b0010010001100000000000000000000000000000000000000000000000000000;
					GGR[3584:3647] <= 64'b0010011000110000000000000000000000000000000000000000000000000000;
					GGR[3648:3711] <= 64'b0010001100001110000000000000000000000000000000000000000000000000;
					GGR[3712:3775] <= 64'b0011000011000000000000000000000000000000000000000000000000000000;
					GGR[3776:3839] <= 64'b0001100000000000000000000000000000000000000000000000000000000000;
					GGR[3840:3903] <= 64'b0000100000000000000000000000000000000000000000000000000000000000;
					GGR[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				1: begin
					GGR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[  64: 127] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[ 128: 191] <= 64'b0000000000000000000000000000011111110000000000000000000000000000;
					GGR[ 192: 255] <= 64'b0000000000000000000000000001110000000000000000000000000000000000;
					GGR[ 256: 319] <= 64'b0000000001111111111000000011000011111100000000000000000000000000;
					GGR[ 320: 383] <= 64'b0000000011000000001100000000001110000100000000000000000000000000;
					GGR[ 384: 447] <= 64'b0000000110000000000100000000000001111111100000000000000000000000;
					GGR[ 448: 511] <= 64'b0000001100000000000110000000000011000000010000000000000000000000;
					GGR[ 512: 575] <= 64'b0000011000000000000010000000000000000000000000000000000000000000;
					GGR[ 576: 639] <= 64'b0000110000000000000110000000000000000000000000000000000000000000;
					GGR[ 640: 703] <= 64'b0000100000000000001100000000000000000000000000000000000000000000;
					GGR[ 704: 767] <= 64'b0001100000000001111000000000000000000000000000000000000000000000;
					GGR[ 768: 831] <= 64'b0001000000000111100001111111111111111111110000000000000000000000;
					GGR[ 832: 895] <= 64'b0001000000001110000011000000011100010000001111000000000000000000;
					GGR[ 896: 959] <= 64'b0001000000110000000110000000000100001100000000111100000000000000;
					GGR[ 960:1023] <= 64'b0011000001100000111100000000000110000100000000000111000000000000;
					GGR[1024:1087] <= 64'b0010000001000011100000000000000011000010000000000001100000000000;
					GGR[1088:1151] <= 64'b0010000011000110000000000000000001100001000000000000111000000000;
					GGR[1152:1215] <= 64'b0010000010011000000000000000000000100000100000000000011100000000;
					GGR[1216:1279] <= 64'b0010000010010000000000000000000000010000100000000000011110000000;
					GGR[1280:1343] <= 64'b0010000011100000000000000000000000011000100000000000001111000000;
					GGR[1344:1407] <= 64'b0011000011100000111100000001111000001000010000000000000101100000;
					GGR[1408:1471] <= 64'b0001000001000001111110000011111100000100010000000000000110110000;
					GGR[1472:1535] <= 64'b0000100001000011111111000011111110000100011000000000000010011000;
					GGR[1536:1599] <= 64'b0000011010000011111111000111111110000100001000000000000011001000;
					GGR[1600:1663] <= 64'b0000001110000010011111000110011110000100001000000000000001000100;
					GGR[1664:1727] <= 64'b0000000110000010011111000110011110000100001000000000000001000100;
					GGR[1728:1791] <= 64'b0000000010000011111111000011111110000100001000000000000001000110;
					GGR[1792:1855] <= 64'b0000000100000001111110000001111100000100001000000000000001000010;
					GGR[1856:1919] <= 64'b0000000100000000000000000000000000000100001000000000000001000010;
					GGR[1920:1983] <= 64'b0000000100000000000000000000000000000100001000000000000001000010;
					GGR[1984:2047] <= 64'b0000000100000110000000110000000001100100001000000000000001000010;
					GGR[2048:2111] <= 64'b0000000100000011000001111000000001000100001000000000000001000010;
					GGR[2112:2175] <= 64'b0000000100000001000011001000000011000100001000000000000001000010;
					GGR[2176:2239] <= 64'b0000000100000001100110001100000110001100001000000000000001000010;
					GGR[2240:2303] <= 64'b0111100010000001111100000111111110001000011000000000000001000010;
					GGR[2304:2367] <= 64'b0100100010000001000000000000000100001000110000000000000001000010;
					GGR[2368:2431] <= 64'b0100010011000001100000000000001100001000100000000000000001000010;
					GGR[2432:2495] <= 64'b1000010001000000100000000000011000011001100000000000000001000110;
					GGR[2496:2559] <= 64'b1000010001000000100000000000110000110001000000000000000011000100;
					GGR[2560:2623] <= 64'b1000001000100000010000000000100000100001000000000000000110001000;
					GGR[2624:2687] <= 64'b1100001110100000011000000011100001100011000000000000001100011000;
					GGR[2688:2751] <= 64'b1100000010010000001111111110000011000010000000000000001000010000;
					GGR[2752:2815] <= 64'b0110000011011000000000000000000010000110000000000000011001100000;
					GGR[2816:2879] <= 64'b0010000001111110000000000000001110001100000000000000010011000000;
					GGR[2880:2943] <= 64'b0010000000011111100000000000010000001000000000000000110110000000;
					GGR[2944:3007] <= 64'b0011000000000001111110000000110000011000000000000001111100000000;
					GGR[3008:3071] <= 64'b0001000000000000000011110001100000110000000000000011110000000000;
					GGR[3072:3135] <= 64'b0001100000000000000001111111111001100000000000000111000000000000;
					GGR[3136:3199] <= 64'b0001111100000000000000000001111111000000000000111100000000000000;
					GGR[3200:3263] <= 64'b0000000111000000000000000111000111111111111111110000000000000000;
					GGR[3264:3327] <= 64'b0000000000111110000001111000000000000000000000000000000000000000;
					GGR[3328:3391] <= 64'b0000000100000011111110000000000000000000000000000000000000000000;
					GGR[3392:3455] <= 64'b0000000100000000000000000000000000000000000000000000000000000000;
					GGR[3456:3519] <= 64'b0010000110000000000000000000000000000000000000000000000000000000;
					GGR[3520:3583] <= 64'b0001110001111000000000000000000000000000000000000000000000000000;
					GGR[3584:3647] <= 64'b0000011100000000000000000000000000000000000000000000000000000000;
					GGR[3648:3711] <= 64'b0000000111000000000000000000000000000000000000000000000000000000;
					GGR[3712:3775] <= 64'b0000000000100000000000000000000000000000000000000000000000000000;
					GGR[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				2: begin
					GGR[   0:  63] <= 64'b0000000000000000000000000000000111111000000000000000000000000000;
					GGR[  64: 127] <= 64'b0000000000000000000000000000011100001110000000000000000000000000;
					GGR[ 128: 191] <= 64'b0000000000000000000000000001100000000010000000000000000000000000;
					GGR[ 192: 255] <= 64'b0000000000000000000000000011000000000010000000000000000000000000;
					GGR[ 256: 319] <= 64'b0000000000000000000000000110000000000110000000000000000000000000;
					GGR[ 320: 383] <= 64'b0000000000000000000000001100000000001100000000000000000000000000;
					GGR[ 384: 447] <= 64'b0000000000000000000000001000000000011000000000000000000000000000;
					GGR[ 448: 511] <= 64'b0000000000000000000000011000000000100000000000000000000000000000;
					GGR[ 512: 575] <= 64'b0000000000000000000000110000000001000000000000000000000000000000;
					GGR[ 576: 639] <= 64'b0000000000000000000001100000000001000000000000000000000000000000;
					GGR[ 640: 703] <= 64'b0000000000000000000001100000000010000000000000000000000000000000;
					GGR[ 704: 767] <= 64'b0000000000000000000001000000000110000000000000000000000000000000;
					GGR[ 768: 831] <= 64'b0000000000000000111111000000000111111111110000000000000000000000;
					GGR[ 832: 895] <= 64'b0000000000000001100001000000000100011000001111000000000000000000;
					GGR[ 896: 959] <= 64'b0000000000000010000001000000001100001100000000111100000000000000;
					GGR[ 960:1023] <= 64'b0000000000001100000001000000001010000100000000000111000000000000;
					GGR[1024:1087] <= 64'b0000000000011000000001000000001011000010000000000001100000000000;
					GGR[1088:1151] <= 64'b0000000001100000000001000000001001100001000000000000111000000000;
					GGR[1152:1215] <= 64'b0000000011000000000001000000001001100000100000000000011100000000;
					GGR[1216:1279] <= 64'b0000000010000000000001000000001000010000100000000000011110000000;
					GGR[1280:1343] <= 64'b0000000110000000000001000000001000011000100000000000001111000000;
					GGR[1344:1407] <= 64'b0000000100000000011111000000001000001000010000000000000101100000;
					GGR[1408:1471] <= 64'b0000001000000001111111000000001000000100010000000000000110110000;
					GGR[1472:1535] <= 64'b0000001000000011111110000000001000000100011000000000000010011000;
					GGR[1536:1599] <= 64'b0000011000000011111111000000001000000100001000000000000011001000;
					GGR[1600:1663] <= 64'b0000010000000010011111000000001000000100001000000000000001000100;
					GGR[1664:1727] <= 64'b0000010000000010011111000000001000000100001000000000000001000100;
					GGR[1728:1791] <= 64'b0000010000000011111110000000001100000100001000000000000001000110;
					GGR[1792:1855] <= 64'b0000010000000001111111000000000100000100001000000000000001000010;
					GGR[1856:1919] <= 64'b0000010000000000000001000000000100000100001000000000000001000010;
					GGR[1920:1983] <= 64'b0000010000000000000001000000000100000100001000000000000001000010;
					GGR[1984:2047] <= 64'b0000010000001000000000100000000010000100001000000000000001000010;
					GGR[2048:2111] <= 64'b0000010000001100000000110000000010000100001000000000000001000010;
					GGR[2112:2175] <= 64'b0000010000000110000011110000000001000100001000000000000001000010;
					GGR[2176:2239] <= 64'b0000010000000111001110011000000000101100001000000000000001000010;
					GGR[2240:2303] <= 64'b0000010000000111111000011000000000111000011000000000000001000010;
					GGR[2304:2367] <= 64'b0000010000000010000000001000000000110000110000000000000001000010;
					GGR[2368:2431] <= 64'b0000010000000010000000001100000000010000100000000000000001000010;
					GGR[2432:2495] <= 64'b0000010000000010000000000100000000011001100000000000000001000010;
					GGR[2496:2559] <= 64'b0000010000000011000000000110000000001001000000000000000011000010;
					GGR[2560:2623] <= 64'b0000011000000001100000000110000000001001000000000000000110000010;
					GGR[2624:2687] <= 64'b0000001000000000110000000110000000001111000000000000001100000110;
					GGR[2688:2751] <= 64'b0000001000000000011111111111000000000010000000000000011000000110;
					GGR[2752:2815] <= 64'b0000001100000000000000000001000000000010000000000000110000011100;
					GGR[2816:2879] <= 64'b0000000110000000000000000001100000000011000000000011100000010000;
					GGR[2880:2943] <= 64'b0000001111000000000000000000110000000001110000000011000001110000;
					GGR[2944:3007] <= 64'b0000011001100000000000000001111000000000001110001110000011000000;
					GGR[3008:3071] <= 64'b0000110000100000000000000111001100000000000011111100001110000000;
					GGR[3072:3135] <= 64'b0011000000111000000000001100000110000000000000000000011000000000;
					GGR[3136:3199] <= 64'b0010000000001100000000001000000011111000000000000000110000000000;
					GGR[3200:3263] <= 64'b0110000001111110000000111000001110001100000000000001100000000000;
					GGR[3264:3327] <= 64'b1100000111000011111111111111111111111111111111111111000000000000;
					GGR[3328:3391] <= 64'b1000000100000000000000000000000000000000000000000000000000000000;
					GGR[3392:3455] <= 64'b1000000100000000000000000000000000000000000000000000000000000000;
					GGR[3456:3519] <= 64'b1000000111000000000000000000000000000000000000000000000000000000;
					GGR[3520:3583] <= 64'b1000000001100000000000000000000000000000000000000000000000000000;
					GGR[3584:3647] <= 64'b1000000000110000000000000000000000000000000000000000000000000000;
					GGR[3648:3711] <= 64'b1000000000011000000000000000000000000000000000000000000000000000;
					GGR[3712:3775] <= 64'b1000000000001000000000000000000000000000000000000000000000000000;
					GGR[3776:3839] <= 64'b1100000000001000000000000000000000000000000000000000000000000000;
					GGR[3840:3903] <= 64'b0111000000011000000000000000000000000000000000000000000000000000;
					GGR[3904:3967] <= 64'b0001111111110000000000000000000000000000000000000000000000000000;
					GGR[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				3: begin
					GGR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[  64: 127] <= 64'b0000000000000000000000000011111000000000000000000000000000000000;
					GGR[ 128: 191] <= 64'b0000000000000000000000111100001110000000000000000000000000000000;
					GGR[ 192: 255] <= 64'b0000000000000000000111000000000010000000000000000000000000000000;
					GGR[ 256: 319] <= 64'b0000000000000000011100000000000001000000000000000000000000000000;
					GGR[ 320: 383] <= 64'b0000000000000000110000000000000001000000000000000000000000000000;
					GGR[ 384: 447] <= 64'b0000000000000000100000000000000011000000000000000000000000000000;
					GGR[ 448: 511] <= 64'b0000000000000001000000011000000010000000000000000000000000000000;
					GGR[ 512: 575] <= 64'b0000000000000010000001111110011110000000000000000000000000000000;
					GGR[ 576: 639] <= 64'b0000000000000110000011000011110000000000000000000000000000000000;
					GGR[ 640: 703] <= 64'b0000000000000100000110000000000000000000000000000000000000000000;
					GGR[ 704: 767] <= 64'b0000000000000100001100000000000000000000000000000000000000000000;
					GGR[ 768: 831] <= 64'b0000000000000100111111111111111111111111110000000000000000000000;
					GGR[ 832: 895] <= 64'b0000000000001101100000000000011100011000001111000000000000000000;
					GGR[ 896: 959] <= 64'b0000000000000110000000000000000100001100000000111100000000000000;
					GGR[ 960:1023] <= 64'b0000000000001100000000000000000110000100000000000111000000000000;
					GGR[1024:1087] <= 64'b0000000000011000000000000000000011000010000000000001100000000000;
					GGR[1088:1151] <= 64'b0000000001100000000000000000000001100001000000000000111000000000;
					GGR[1152:1215] <= 64'b0000000011000000000000000000000001100000100000000000011100000000;
					GGR[1216:1279] <= 64'b0000000010000000000000000000000000010000100000000000011110000000;
					GGR[1280:1343] <= 64'b0000000110000000000000000000000000011000100000000000001111000000;
					GGR[1344:1407] <= 64'b0000000100000000011100000001111000001000010000000000000101100000;
					GGR[1408:1471] <= 64'b0000001000000001111110000011111100000100010000000000000110110000;
					GGR[1472:1535] <= 64'b0000001000000011111110000011111110000100011000000000000010011000;
					GGR[1536:1599] <= 64'b0000011000000011111111000111111110000100001000000000000011001000;
					GGR[1600:1663] <= 64'b0000010000000010011111000110011110000100001000000000000001000100;
					GGR[1664:1727] <= 64'b0000010000000010011111000110011110000100001000000000000001000100;
					GGR[1728:1791] <= 64'b0000010000000011111110000011111110000100001000000000000001000110;
					GGR[1792:1855] <= 64'b0000010000000001111110000001111100000100001000000000000001000010;
					GGR[1856:1919] <= 64'b0000010000000000000000000000000000100100001000000000000001000010;
					GGR[1920:1983] <= 64'b0000010000000000000000000000000001100100001000000000000001000010;
					GGR[1984:2047] <= 64'b0000010000001000000000000000000011000100001000000000000001000010;
					GGR[2048:2111] <= 64'b0000010000001100000000000000000110000100001000000000000001000010;
					GGR[2112:2175] <= 64'b0000010000000110000011111000011100000100001000000000000001000010;
					GGR[2176:2239] <= 64'b0000010000000111001110001100110100001100001000000000000001000010;
					GGR[2240:2303] <= 64'b0000010000000111111000000111100100001000011000000000000001000010;
					GGR[2304:2367] <= 64'b0000010000000010000000000000001100001000110000000000000001000010;
					GGR[2368:2431] <= 64'b0000010000000010000000000000001000001000100000000000000001000010;
					GGR[2432:2495] <= 64'b0000010000000010000000000000011000011001100000000000000001000010;
					GGR[2496:2559] <= 64'b0000010000000011000000000000110000110001000000000000000011000010;
					GGR[2560:2623] <= 64'b0000011000000001100000000001100000100001000000000000000110000010;
					GGR[2624:2687] <= 64'b0000001000000000110000000111000001100011000000000000001100000110;
					GGR[2688:2751] <= 64'b0000001000000000011111111100000011000010000000000000011000000110;
					GGR[2752:2815] <= 64'b0000001100000000000000000000000010000110000000000000110000011100;
					GGR[2816:2879] <= 64'b0000000110000000000000000000001110001100000000000011100000010000;
					GGR[2880:2943] <= 64'b0000000011000000000000000000011100001000000000000011000001110000;
					GGR[2944:3007] <= 64'b0000000001100000000000000001111000011000000000001110000011000000;
					GGR[3008:3071] <= 64'b0000000000100000000000000011100000110000000000011100001110000000;
					GGR[3072:3135] <= 64'b0000000000111000000000000110000001100000000001110000011000000000;
					GGR[3136:3199] <= 64'b0000000000001100000000001000000111000000000111000000110000000000;
					GGR[3200:3263] <= 64'b0001111110000110000000011000000100000000001100000001100000000000;
					GGR[3264:3327] <= 64'b0011000010000011111111100000001111111111111111111111000000000000;
					GGR[3328:3391] <= 64'b0110000010000000000001100000011000000000000000000000000000000000;
					GGR[3392:3455] <= 64'b0100000110000000000110000000110000000000000000000000000000000000;
					GGR[3456:3519] <= 64'b1000000100000000001100000001100000000000000000000000000000000000;
					GGR[3520:3583] <= 64'b1000000111100000011000000011000000000000000000000000000000000000;
					GGR[3584:3647] <= 64'b1000000001111111100000000010000000000000000000000000000000000000;
					GGR[3648:3711] <= 64'b1100000000000000000000000110000000000000000000000000000000000000;
					GGR[3712:3775] <= 64'b0100000000000000000000001100000000000000000000000000000000000000;
					GGR[3776:3839] <= 64'b0110000000000000000000110000000000000000000000000000000000000000;
					GGR[3840:3903] <= 64'b0011100000000000000011100000000000000000000000000000000000000000;
					GGR[3904:3967] <= 64'b0000111100000000011110000000000000000000000000000000000000000000;
					GGR[3968:4031] <= 64'b0000000111111111100000000000000000000000000000000000000000000000;
					GGR[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				4: begin
					GGR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[  64: 127] <= 64'b0000000000000111111000000000000000000000000000000000000000000000;
					GGR[ 128: 191] <= 64'b0000000001111000001100000000000000000000000000000000000000000000;
					GGR[ 192: 255] <= 64'b0000000111000000001100000000000000000000000000000000000000000000;
					GGR[ 256: 319] <= 64'b0000001100000000011000000000000000000000000000000000000000000000;
					GGR[ 320: 383] <= 64'b0000110000000000110000000000000000000000000000000000000000000000;
					GGR[ 384: 447] <= 64'b0000100000000000100000000000000000000000000000000000000000000000;
					GGR[ 448: 511] <= 64'b0000100000000001000000000000000000000000000000000000000000000000;
					GGR[ 512: 575] <= 64'b0001000000000011000000000000000000000000000000000000000000000000;
					GGR[ 576: 639] <= 64'b0001000000000110000000000000000000000000000000000000000000000000;
					GGR[ 640: 703] <= 64'b0001000000000100000000000000000000000000000000000000000000000000;
					GGR[ 704: 767] <= 64'b0001000000000100000000000000000000000000000000000000000000000000;
					GGR[ 768: 831] <= 64'b0001000000000100000001111111111111111111110000000000000000000000;
					GGR[ 832: 895] <= 64'b0011000000000100000011000000011100010000001111000000000000000000;
					GGR[ 896: 959] <= 64'b0010000000001100000110000000000100001100000000111100000000000000;
					GGR[ 960:1023] <= 64'b0010000000001000111100000000000110000100000000000111000000000000;
					GGR[1024:1087] <= 64'b0010000000001011100000000000000011000010000000000001100000000000;
					GGR[1088:1151] <= 64'b0010000000001110000000000000000001100001000000000000111000000000;
					GGR[1152:1215] <= 64'b0010000000011000000000000000000000100000100000000000011100000000;
					GGR[1216:1279] <= 64'b0010000000010000000000000000000000010000100000000000011110000000;
					GGR[1280:1343] <= 64'b0010000000010000000000000000000000011000100000000000001111000000;
					GGR[1344:1407] <= 64'b0010000000010000111100000001111000001000010000000000000101100000;
					GGR[1408:1471] <= 64'b0010000000010001111110000011111100000100010000000000000110110000;
					GGR[1472:1535] <= 64'b0010000000010011111111000011111110000100011000000000000010011000;
					GGR[1536:1599] <= 64'b0010000000010011111111000111111110000100001000000000000011001000;
					GGR[1600:1663] <= 64'b0010000000010010011111000110011110000100001000000000000001000100;
					GGR[1664:1727] <= 64'b0010000000010010011111000110011110000100001000000000000001000100;
					GGR[1728:1791] <= 64'b0011000000010011111111000011111110000100001000000000000001000110;
					GGR[1792:1855] <= 64'b0001000000010001111110000001111100000100001000000000000001000010;
					GGR[1856:1919] <= 64'b0001000000010000000000000000000000000100001000000000000001000010;
					GGR[1920:1983] <= 64'b0001000000011010000000000000000000000100001000000000000001000010;
					GGR[1984:2047] <= 64'b0001000000001011000000110000000001100100001000000000000001000010;
					GGR[2048:2111] <= 64'b0001000000001101100011111110000001000100001000000000000001000010;
					GGR[2112:2175] <= 64'b0000100000000100111110000011000011000100001000000000000001000010;
					GGR[2176:2239] <= 64'b0000100000000110100000000001111110001100001000000000000001000010;
					GGR[2240:2303] <= 64'b0000110000000010110000000000000110001000011000000000000001000010;
					GGR[2304:2367] <= 64'b0000010000000001010000000000000100001000110000000000000001000010;
					GGR[2368:2431] <= 64'b0000011000000001101000000000001100001000100000000000000001000010;
					GGR[2432:2495] <= 64'b0000001000000000110110000000011000011001100000000000000001000010;
					GGR[2496:2559] <= 64'b0000001100000000011011000000110000110001000000000000000011000010;
					GGR[2560:2623] <= 64'b0000000100000000001101111111100000100001000000000000000110000010;
					GGR[2624:2687] <= 64'b0000000100000000000110000000000001100011000000000000001100000110;
					GGR[2688:2751] <= 64'b0011110011000000000011100000000011000010000000000000001000000110;
					GGR[2752:2815] <= 64'b0110011001110000000001100000000010000110000000000000011000011100;
					GGR[2816:2879] <= 64'b0100001100011000000000110000001110001100000000000000010000011000;
					GGR[2880:2943] <= 64'b1000000110001110000000011100010000001000000000000001110000110000;
					GGR[2944:3007] <= 64'b1000000011000011100000000111110000011000000000000011000001110000;
					GGR[3008:3071] <= 64'b1000000001100000111100000001100000110000000000000110000011100000;
					GGR[3072:3135] <= 64'b1000000000111100000110000000111001100000000000001100000011000000;
					GGR[3136:3199] <= 64'b1000000000000111000011000000000111000000000001111100001110000000;
					GGR[3200:3263] <= 64'b0110000000000000111111111111111111111111111111110000011100000000;
					GGR[3264:3327] <= 64'b0110000000000000000000000000000000000000000000000011111000000000;
					GGR[3328:3391] <= 64'b0011100000000000000000000000000000000000000000000111100000000000;
					GGR[3392:3455] <= 64'b0000111000000000000000000000000000000000000000111100000000000000;
					GGR[3456:3519] <= 64'b0000001111000000000000000000000000000000011111100000000000000000;
					GGR[3520:3583] <= 64'b0000000011000000000000000000000000000001111000000000000000000000;
					GGR[3584:3647] <= 64'b0000000001111000000000000000000001111111000000000000000000000000;
					GGR[3648:3711] <= 64'b0000000000001111111111111111111111000000000000000000000000000000;
					GGR[3712:3775] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3776:3839] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3840:3903] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3904:3967] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[3968:4031] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[4032:4095] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
				end
				default: begin
					GGR[   0:  63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
					GGR[  64: 127] <= 64'b0000000000000000000000000010010001100111111110000000000000000000;
					GGR[ 128: 191] <= 64'b0000000000000000000000001110110010001100000011000000000000000000;
					GGR[ 192: 255] <= 64'b0000000000000000000000001001100100011000000001000000000000000000;
					GGR[ 256: 319] <= 64'b0000000000000000000000010001001000010000000011000000000000000000;
					GGR[ 320: 383] <= 64'b0000000000000000000000110011001000110000000110000000000000000000;
					GGR[ 384: 447] <= 64'b0000000000000000000000100010011001100000000100000000000000000000;
					GGR[ 448: 511] <= 64'b0000000000000000000001100010010001000000001100000000000000000000;
					GGR[ 512: 575] <= 64'b0000000000000000000000000000000001000000001000000000000000000000;
					GGR[ 576: 639] <= 64'b0000000000000000000000000000000011000000011000000000000000000000;
					GGR[ 640: 703] <= 64'b0000000000000000000000000000000010000000010000000000000000000000;
					GGR[ 704: 767] <= 64'b0000000000000000000000111111111110000000110000000000000000000000;
					GGR[ 768: 831] <= 64'b0000000000000000111111100000011110000000110000000000000000000000;
					GGR[ 832: 895] <= 64'b0000000000000001100000000000001010000000101111000000000000000000;
					GGR[ 896: 959] <= 64'b0000000000000010000000000000001010000000100000111100000000000000;
					GGR[ 960:1023] <= 64'b0000000000001100000000000000000110000000100000000111000000000000;
					GGR[1024:1087] <= 64'b0000000000011000000000000000000010000000100000000001100000000000;
					GGR[1088:1151] <= 64'b0000000001100000000000000000000010000000100000000000111000000000;
					GGR[1152:1215] <= 64'b0000000011000000000000000000000110000000100000000000011100000000;
					GGR[1216:1279] <= 64'b0000000010000000000000000000000100000000110000000000011110000000;
					GGR[1280:1343] <= 64'b0000000110000011100000000111000100000000110000000000001111000000;
					GGR[1344:1407] <= 64'b0000000100001111111000001111110100000000010000000000000101100000;
					GGR[1408:1471] <= 64'b0000001000011111111000011111111100000000010000000000000110110000;
					GGR[1472:1535] <= 64'b0000001000011111111100011111111100000000011000000000000010011000;
					GGR[1536:1599] <= 64'b0000011000111111111100111111111100000000001000000000000011001100;
					GGR[1600:1663] <= 64'b0000010000111001111100111001111100000000001000000000000001000100;
					GGR[1664:1727] <= 64'b0000010000111001111100111001111110000000001000000000000001000100;
					GGR[1728:1791] <= 64'b0000010000011111111100011111111110000000001000000000000001000110;
					GGR[1792:1855] <= 64'b0000010000011111111000011111111110000000001100000000000001000010;
					GGR[1856:1919] <= 64'b0000010000000011111000000011111001000000000110000000000001000010;
					GGR[1920:1983] <= 64'b0000010000000000000000000000000001000000000010000000000001000010;
					GGR[1984:2047] <= 64'b0000010000001000000000000000000101000000000010000000000001000010;
					GGR[2048:2111] <= 64'b0000010000001000000001100000001100100000000010000000000001000010;
					GGR[2112:2175] <= 64'b0000010000000100000011110000001100100000000010000000000001000010;
					GGR[2176:2239] <= 64'b0000010000000110001110011000111000100000000011000000000001000010;
					GGR[2240:2303] <= 64'b0000010000000111111000001111111000010000000001000000000001000010;
					GGR[2304:2367] <= 64'b0000010000000010000000000000010000010000000001000000000001000010;
					GGR[2368:2431] <= 64'b0000010000000010000000000000010000011000000001100000000001000010;
					GGR[2432:2495] <= 64'b0000010000000010000000000000110000011000000000110000000001000010;
					GGR[2496:2559] <= 64'b0000010000000011000000000001100000010100000000010000000011000010;
					GGR[2560:2623] <= 64'b0000011000000001100000000011000000001111000000011000000110000010;
					GGR[2624:2687] <= 64'b0000001000000000110000000110000000011011000000001100000100000010;
					GGR[2688:2751] <= 64'b0000001000000000011111111000000000110011100000000110011100000010;
					GGR[2752:2815] <= 64'b0000001100000000000000000000000001100010110000000011111000000110;
					GGR[2816:2879] <= 64'b0000000110000000000000000000000011000110011000000000110000000100;
					GGR[2880:2943] <= 64'b0000000011000000000000000000000010000100001100000001100000011100;
					GGR[2944:3007] <= 64'b0000000001100000000000000000001100011000000110000110000000011000;
					GGR[3008:3071] <= 64'b0000000000100000000000000000001000010000000011001100000000110000;
					GGR[3072:3135] <= 64'b0000000001111000000000000000110001110000000001111000000001100000;
					GGR[3136:3199] <= 64'b0000000000001100000000000001100011000000000000110000000110000000;
					GGR[3200:3263] <= 64'b0000000010000010000000000110000110000000000011100000011100000000;
					GGR[3264:3327] <= 64'b0000001000000011111111111111111111111111111111111111110000000000;
					GGR[3328:3391] <= 64'b0000001000000000110000000000000000000000000000000000000000000000;
					GGR[3392:3455] <= 64'b0000010000000000100000000000000000000000000000000000000000000000;
					GGR[3456:3519] <= 64'b0000010000000000110000000000000000000000000000000000000000000000;
					GGR[3520:3583] <= 64'b0000010000000000010000000000000000000000000000000000000000000000;
					GGR[3584:3647] <= 64'b0000010000000000011100000000000000000000000000000000000000000000;
					GGR[3648:3711] <= 64'b0000010000000000000111100000000000000000000000000000000000000000;
					GGR[3712:3775] <= 64'b0000110000000000000000111000000000000000000000000000000000000000;
					GGR[3776:3839] <= 64'b0000001000000000000000001100000000000000000000000000000000000000;
					GGR[3840:3903] <= 64'b0000001100000000000000000100000000000000000000000000000000000000;
					GGR[3904:3967] <= 64'b0000000111000000000000001100000000000000000000000000000000000000;
					GGR[3968:4031] <= 64'b0000000000111000000000011000000000000000000000000000000000000000;
					GGR[4032:4095] <= 64'b0000000000000111111111100000000000000000000000000000000000000000;
				end
			endcase
		end
		else begin
		end
		if(count==3'b110)
			count <= 3'b000;
		else
			count <= (count+1);
		if(display==10)
			display <= 0;
		else 
			display <= (display+1);
	end
	
	
endmodule
